magic
tech sky130A
timestamp 1699645850
<< nwell >>
rect -110 135 295 275
<< nmos >>
rect 0 -15 15 85
rect 145 -15 160 85
rect 210 -15 225 85
<< pmos >>
rect 0 155 15 255
rect 145 155 160 255
rect 210 155 225 255
<< ndiff >>
rect -50 70 0 85
rect -50 0 -35 70
rect -15 0 0 70
rect -50 -15 0 0
rect 15 70 60 85
rect 100 70 145 85
rect 15 0 30 70
rect 50 0 60 70
rect 100 0 110 70
rect 130 0 145 70
rect 15 -15 60 0
rect 100 -15 145 0
rect 160 70 210 85
rect 160 0 175 70
rect 195 0 210 70
rect 160 -15 210 0
rect 225 70 275 85
rect 225 0 240 70
rect 260 0 275 70
rect 225 -15 275 0
<< pdiff >>
rect -45 240 0 255
rect -45 170 -35 240
rect -15 170 0 240
rect -45 155 0 170
rect 15 240 65 255
rect 15 170 30 240
rect 50 170 65 240
rect 15 155 65 170
rect 95 240 145 255
rect 95 170 110 240
rect 130 170 145 240
rect 95 155 145 170
rect 160 240 210 255
rect 160 170 175 240
rect 195 170 210 240
rect 160 155 210 170
rect 225 240 275 255
rect 225 170 240 240
rect 260 170 275 240
rect 225 155 275 170
<< ndiffc >>
rect -35 0 -15 70
rect 30 0 50 70
rect 110 0 130 70
rect 175 0 195 70
rect 240 0 260 70
<< pdiffc >>
rect -35 170 -15 240
rect 30 170 50 240
rect 110 170 130 240
rect 175 170 195 240
rect 240 170 260 240
<< psubdiff >>
rect 60 70 100 85
rect 60 0 70 70
rect 90 0 100 70
rect 60 -15 100 0
<< nsubdiff >>
rect -90 240 -45 255
rect -90 170 -75 240
rect -55 170 -45 240
rect -90 155 -45 170
<< psubdiffcont >>
rect 70 0 90 70
<< nsubdiffcont >>
rect -75 170 -55 240
<< poly >>
rect 0 295 225 310
rect 0 255 15 295
rect 145 255 160 270
rect 210 255 225 295
rect 0 85 15 155
rect 145 135 160 155
rect 60 130 160 135
rect 60 110 70 130
rect 90 110 160 130
rect 60 105 160 110
rect 145 85 160 105
rect 210 85 225 155
rect 0 -30 15 -15
rect 145 -30 160 -15
rect 210 -30 225 -15
<< polycont >>
rect 70 110 90 130
<< locali >>
rect -85 240 -5 250
rect -85 170 -75 240
rect -55 170 -35 240
rect -15 170 -5 240
rect -85 160 -5 170
rect 20 240 60 250
rect 20 170 30 240
rect 50 170 60 240
rect 20 160 60 170
rect 100 240 140 250
rect 100 170 110 240
rect 130 170 140 240
rect 100 160 140 170
rect 165 240 205 250
rect 165 170 175 240
rect 195 170 205 240
rect 40 135 60 160
rect -25 130 100 135
rect -25 110 70 130
rect 90 110 100 130
rect -25 105 100 110
rect -25 80 -5 105
rect -45 70 -5 80
rect -45 0 -35 70
rect -15 0 -5 70
rect -45 -10 -5 0
rect 20 70 140 80
rect 20 0 30 70
rect 50 0 70 70
rect 90 0 110 70
rect 130 0 140 70
rect 20 -10 140 0
rect 165 70 205 170
rect 230 240 270 250
rect 230 170 240 240
rect 260 170 270 240
rect 230 160 270 170
rect 165 0 175 70
rect 195 0 205 70
rect 165 -10 205 0
rect 230 70 270 80
rect 230 0 240 70
rect 260 0 270 70
rect 230 -10 270 0
<< viali >>
rect -75 170 -55 240
rect -35 170 -15 240
rect 110 170 130 240
rect 30 0 50 70
rect 70 0 90 70
rect 110 0 130 70
rect 240 170 260 240
rect 240 0 260 70
<< metal1 >>
rect -85 245 -5 250
rect -85 165 -80 245
rect -50 165 -40 245
rect -10 165 -5 245
rect -85 160 -5 165
rect 100 240 140 250
rect 100 170 110 240
rect 130 170 140 240
rect 100 160 140 170
rect 230 245 270 250
rect 230 165 235 245
rect 265 165 270 245
rect 230 160 270 165
rect 120 135 140 160
rect 120 115 250 135
rect 230 80 250 115
rect 15 75 145 80
rect 15 -5 20 75
rect 50 -5 65 75
rect 95 -5 110 75
rect 140 -5 145 75
rect 15 -10 145 -5
rect 230 70 270 80
rect 230 0 240 70
rect 260 0 270 70
rect 230 -10 270 0
<< via1 >>
rect -80 240 -50 245
rect -80 170 -75 240
rect -75 170 -55 240
rect -55 170 -50 240
rect -80 165 -50 170
rect -40 240 -10 245
rect -40 170 -35 240
rect -35 170 -15 240
rect -15 170 -10 240
rect -40 165 -10 170
rect 235 240 265 245
rect 235 170 240 240
rect 240 170 260 240
rect 260 170 265 240
rect 235 165 265 170
rect 20 70 50 75
rect 20 0 30 70
rect 30 0 50 70
rect 20 -5 50 0
rect 65 70 95 75
rect 65 0 70 70
rect 70 0 90 70
rect 90 0 95 70
rect 65 -5 95 0
rect 110 70 140 75
rect 110 0 130 70
rect 130 0 140 70
rect 110 -5 140 0
<< metal2 >>
rect -85 245 -5 250
rect -85 165 -80 245
rect -50 165 -40 245
rect -10 165 -5 245
rect -85 160 -5 165
rect 230 245 270 250
rect 230 165 235 245
rect 265 165 270 245
rect 230 160 270 165
rect 230 115 250 160
rect 125 95 250 115
rect 125 80 145 95
rect 15 75 145 80
rect 15 -5 20 75
rect 50 -5 65 75
rect 95 -5 110 75
rect 140 -5 145 75
rect 15 -10 145 -5
<< labels >>
rlabel locali 185 250 185 250 1 Y
port 1 n
rlabel metal1 270 35 270 35 3 Vbn
port 2 e
rlabel poly 5 -30 5 -30 5 S
port 3 s
rlabel metal2 -85 205 -85 205 7 VP
port 4 w
rlabel metal2 145 35 145 35 3 VN
port 5 e
<< end >>
