magic
tech sky130A
timestamp 1699582308
<< nmos >>
rect -155 0 -55 1200
rect -5 0 95 1200
rect 145 0 245 1200
rect 295 0 395 1200
rect 445 0 545 1200
rect 675 0 775 1200
rect 825 0 925 1200
rect 975 0 1075 1200
rect 1125 0 1225 1200
rect 1405 0 1505 1200
rect 1555 0 1655 1200
rect 1705 0 1805 1200
rect 1855 0 1955 1200
rect 2005 0 2105 1200
rect 2155 0 2255 1200
rect 2305 0 2405 1200
rect 2455 0 2555 1200
rect 2605 0 2705 1200
rect 2755 0 2855 1200
rect 2905 0 3005 1200
rect 3055 0 3155 1200
rect 3205 0 3305 1200
rect 3355 0 3455 1200
rect 3505 0 3605 1200
rect 3655 0 3755 1200
rect 3805 0 3905 1200
rect 3955 0 4055 1200
rect 4205 0 4305 1200
rect 4355 0 4455 1200
rect 4505 0 4605 1200
rect 4655 0 4755 1200
rect 4805 0 4905 1200
rect 4955 0 5055 1200
rect 5105 0 5205 1200
rect -155 -1510 -55 -310
rect -5 -1510 95 -310
rect 225 -1510 325 -310
rect 375 -1510 475 -310
rect 525 -1510 625 -310
rect 675 -1510 775 -310
rect 825 -1510 925 -310
rect 975 -1510 1075 -310
rect 1125 -1510 1225 -310
rect 1275 -1510 1375 -310
rect 1425 -1510 1525 -310
rect 1575 -1510 1675 -310
rect 1725 -1510 1825 -310
rect 1875 -1510 1975 -310
rect 2025 -1510 2125 -310
rect 2175 -1510 2275 -310
rect 2325 -1510 2425 -310
rect 2475 -1510 2575 -310
rect 2755 -1510 2855 -310
rect 2985 -1510 3085 -310
rect 3135 -1510 3235 -310
rect 3285 -1510 3385 -310
rect 3435 -1510 3535 -310
rect 3665 -1510 3765 -310
rect 3815 -1510 3915 -310
rect 3965 -1510 4065 -310
rect 4115 -1510 4215 -310
rect 4265 -1510 4365 -310
rect 4415 -1510 4515 -310
rect 4565 -1510 4665 -310
rect 4715 -1510 4815 -310
rect 4865 -1510 4965 -310
<< ndiff >>
rect -205 1185 -155 1200
rect -205 15 -190 1185
rect -170 15 -155 1185
rect -205 0 -155 15
rect -55 1185 -5 1200
rect -55 15 -40 1185
rect -20 15 -5 1185
rect -55 0 -5 15
rect 95 1185 145 1200
rect 95 15 110 1185
rect 130 15 145 1185
rect 95 0 145 15
rect 245 1185 295 1200
rect 245 15 260 1185
rect 280 15 295 1185
rect 245 0 295 15
rect 395 1185 445 1200
rect 395 15 410 1185
rect 430 15 445 1185
rect 395 0 445 15
rect 545 1185 595 1200
rect 545 15 560 1185
rect 580 15 595 1185
rect 545 0 595 15
rect 625 1185 675 1200
rect 625 15 640 1185
rect 660 15 675 1185
rect 625 0 675 15
rect 775 1185 825 1200
rect 775 15 790 1185
rect 810 15 825 1185
rect 775 0 825 15
rect 925 1185 975 1200
rect 925 15 940 1185
rect 960 15 975 1185
rect 925 0 975 15
rect 1075 1185 1125 1200
rect 1075 15 1090 1185
rect 1110 15 1125 1185
rect 1075 0 1125 15
rect 1225 1185 1275 1200
rect 1225 15 1240 1185
rect 1260 15 1275 1185
rect 1225 0 1275 15
rect 1355 1185 1405 1200
rect 1355 15 1370 1185
rect 1390 15 1405 1185
rect 1355 0 1405 15
rect 1505 1185 1555 1200
rect 1505 15 1520 1185
rect 1540 15 1555 1185
rect 1505 0 1555 15
rect 1655 1185 1705 1200
rect 1655 15 1670 1185
rect 1690 15 1705 1185
rect 1655 0 1705 15
rect 1805 1185 1855 1200
rect 1805 15 1820 1185
rect 1840 15 1855 1185
rect 1805 0 1855 15
rect 1955 1185 2005 1200
rect 1955 15 1970 1185
rect 1990 15 2005 1185
rect 1955 0 2005 15
rect 2105 1185 2155 1200
rect 2105 15 2120 1185
rect 2140 15 2155 1185
rect 2105 0 2155 15
rect 2255 1185 2305 1200
rect 2255 15 2270 1185
rect 2290 15 2305 1185
rect 2255 0 2305 15
rect 2405 1185 2455 1200
rect 2405 15 2420 1185
rect 2440 15 2455 1185
rect 2405 0 2455 15
rect 2555 1185 2605 1200
rect 2555 15 2570 1185
rect 2590 15 2605 1185
rect 2555 0 2605 15
rect 2705 1185 2755 1200
rect 2705 15 2720 1185
rect 2740 15 2755 1185
rect 2705 0 2755 15
rect 2855 1185 2905 1200
rect 2855 15 2870 1185
rect 2890 15 2905 1185
rect 2855 0 2905 15
rect 3005 1185 3055 1200
rect 3005 15 3020 1185
rect 3040 15 3055 1185
rect 3005 0 3055 15
rect 3155 1185 3205 1200
rect 3155 15 3170 1185
rect 3190 15 3205 1185
rect 3155 0 3205 15
rect 3305 1185 3355 1200
rect 3305 15 3320 1185
rect 3340 15 3355 1185
rect 3305 0 3355 15
rect 3455 1185 3505 1200
rect 3455 15 3470 1185
rect 3490 15 3505 1185
rect 3455 0 3505 15
rect 3605 1185 3655 1200
rect 3605 15 3620 1185
rect 3640 15 3655 1185
rect 3605 0 3655 15
rect 3755 1185 3805 1200
rect 3755 15 3770 1185
rect 3790 15 3805 1185
rect 3755 0 3805 15
rect 3905 1185 3955 1200
rect 3905 15 3920 1185
rect 3940 15 3955 1185
rect 3905 0 3955 15
rect 4055 1185 4105 1200
rect 4155 1185 4205 1200
rect 4055 15 4070 1185
rect 4090 15 4105 1185
rect 4155 15 4170 1185
rect 4190 15 4205 1185
rect 4055 0 4105 15
rect 4155 0 4205 15
rect 4305 1185 4355 1200
rect 4305 15 4320 1185
rect 4340 15 4355 1185
rect 4305 0 4355 15
rect 4455 1185 4505 1200
rect 4455 15 4470 1185
rect 4490 15 4505 1185
rect 4455 0 4505 15
rect 4605 1185 4655 1200
rect 4605 15 4620 1185
rect 4640 15 4655 1185
rect 4605 0 4655 15
rect 4755 1185 4805 1200
rect 4755 15 4770 1185
rect 4790 15 4805 1185
rect 4755 0 4805 15
rect 4905 1185 4955 1200
rect 4905 15 4920 1185
rect 4940 15 4955 1185
rect 4905 0 4955 15
rect 5055 1185 5105 1200
rect 5055 15 5070 1185
rect 5090 15 5105 1185
rect 5055 0 5105 15
rect 5205 1185 5255 1200
rect 5205 15 5220 1185
rect 5240 15 5255 1185
rect 5205 0 5255 15
rect -205 -325 -155 -310
rect -205 -1495 -190 -325
rect -170 -1495 -155 -325
rect -205 -1510 -155 -1495
rect -55 -325 -5 -310
rect -55 -1495 -40 -325
rect -20 -1495 -5 -325
rect -55 -1510 -5 -1495
rect 95 -325 145 -310
rect 95 -1495 110 -325
rect 130 -1495 145 -325
rect 95 -1510 145 -1495
rect 175 -325 225 -310
rect 175 -1495 190 -325
rect 210 -1495 225 -325
rect 175 -1510 225 -1495
rect 325 -325 375 -310
rect 325 -1495 340 -325
rect 360 -1495 375 -325
rect 325 -1510 375 -1495
rect 475 -325 525 -310
rect 475 -1495 490 -325
rect 510 -1495 525 -325
rect 475 -1510 525 -1495
rect 625 -325 675 -310
rect 625 -1495 640 -325
rect 660 -1495 675 -325
rect 625 -1510 675 -1495
rect 775 -325 825 -310
rect 775 -1495 790 -325
rect 810 -1495 825 -325
rect 775 -1510 825 -1495
rect 925 -325 975 -310
rect 925 -1495 940 -325
rect 960 -1495 975 -325
rect 925 -1510 975 -1495
rect 1075 -325 1125 -310
rect 1075 -1495 1090 -325
rect 1110 -1495 1125 -325
rect 1075 -1510 1125 -1495
rect 1225 -325 1275 -310
rect 1225 -1495 1240 -325
rect 1260 -1495 1275 -325
rect 1225 -1510 1275 -1495
rect 1375 -325 1425 -310
rect 1375 -1495 1390 -325
rect 1410 -1495 1425 -325
rect 1375 -1510 1425 -1495
rect 1525 -325 1575 -310
rect 1525 -1495 1540 -325
rect 1560 -1495 1575 -325
rect 1525 -1510 1575 -1495
rect 1675 -325 1725 -310
rect 1675 -1495 1690 -325
rect 1710 -1495 1725 -325
rect 1675 -1510 1725 -1495
rect 1825 -325 1875 -310
rect 1825 -1495 1840 -325
rect 1860 -1495 1875 -325
rect 1825 -1510 1875 -1495
rect 1975 -325 2025 -310
rect 1975 -1495 1990 -325
rect 2010 -1495 2025 -325
rect 1975 -1510 2025 -1495
rect 2125 -325 2175 -310
rect 2125 -1495 2140 -325
rect 2160 -1495 2175 -325
rect 2125 -1510 2175 -1495
rect 2275 -325 2325 -310
rect 2275 -1495 2290 -325
rect 2310 -1495 2325 -325
rect 2275 -1510 2325 -1495
rect 2425 -325 2475 -310
rect 2425 -1495 2440 -325
rect 2460 -1495 2475 -325
rect 2425 -1510 2475 -1495
rect 2575 -325 2625 -310
rect 2575 -1495 2590 -325
rect 2610 -1495 2625 -325
rect 2575 -1510 2625 -1495
rect 2705 -325 2755 -310
rect 2705 -1495 2720 -325
rect 2740 -1495 2755 -325
rect 2705 -1510 2755 -1495
rect 2855 -325 2905 -310
rect 2855 -1495 2870 -325
rect 2890 -1495 2905 -325
rect 2855 -1510 2905 -1495
rect 2935 -325 2985 -310
rect 2935 -1495 2950 -325
rect 2970 -1495 2985 -325
rect 2935 -1510 2985 -1495
rect 3085 -325 3135 -310
rect 3085 -1495 3100 -325
rect 3120 -1495 3135 -325
rect 3085 -1510 3135 -1495
rect 3235 -325 3285 -310
rect 3235 -1495 3250 -325
rect 3270 -1495 3285 -325
rect 3235 -1510 3285 -1495
rect 3385 -325 3435 -310
rect 3385 -1495 3400 -325
rect 3420 -1495 3435 -325
rect 3385 -1510 3435 -1495
rect 3535 -325 3585 -310
rect 3535 -1495 3550 -325
rect 3570 -1495 3585 -325
rect 3535 -1510 3585 -1495
rect 3615 -325 3665 -310
rect 3615 -1495 3630 -325
rect 3650 -1495 3665 -325
rect 3615 -1510 3665 -1495
rect 3765 -325 3815 -310
rect 3765 -1495 3780 -325
rect 3800 -1495 3815 -325
rect 3765 -1510 3815 -1495
rect 3915 -325 3965 -310
rect 3915 -1495 3930 -325
rect 3950 -1495 3965 -325
rect 3915 -1510 3965 -1495
rect 4065 -325 4115 -310
rect 4065 -1495 4080 -325
rect 4100 -1495 4115 -325
rect 4065 -1510 4115 -1495
rect 4215 -325 4265 -310
rect 4215 -1495 4230 -325
rect 4250 -1495 4265 -325
rect 4215 -1510 4265 -1495
rect 4365 -325 4415 -310
rect 4365 -1495 4380 -325
rect 4400 -1495 4415 -325
rect 4365 -1510 4415 -1495
rect 4515 -325 4565 -310
rect 4515 -1495 4530 -325
rect 4550 -1495 4565 -325
rect 4515 -1510 4565 -1495
rect 4665 -325 4715 -310
rect 4665 -1495 4680 -325
rect 4700 -1495 4715 -325
rect 4665 -1510 4715 -1495
rect 4815 -325 4865 -310
rect 4815 -1495 4830 -325
rect 4850 -1495 4865 -325
rect 4815 -1510 4865 -1495
rect 4965 -325 5015 -310
rect 4965 -1495 4980 -325
rect 5000 -1495 5015 -325
rect 4965 -1510 5015 -1495
<< ndiffc >>
rect -190 15 -170 1185
rect -40 15 -20 1185
rect 110 15 130 1185
rect 260 15 280 1185
rect 410 15 430 1185
rect 560 15 580 1185
rect 640 15 660 1185
rect 790 15 810 1185
rect 940 15 960 1185
rect 1090 15 1110 1185
rect 1240 15 1260 1185
rect 1370 15 1390 1185
rect 1520 15 1540 1185
rect 1670 15 1690 1185
rect 1820 15 1840 1185
rect 1970 15 1990 1185
rect 2120 15 2140 1185
rect 2270 15 2290 1185
rect 2420 15 2440 1185
rect 2570 15 2590 1185
rect 2720 15 2740 1185
rect 2870 15 2890 1185
rect 3020 15 3040 1185
rect 3170 15 3190 1185
rect 3320 15 3340 1185
rect 3470 15 3490 1185
rect 3620 15 3640 1185
rect 3770 15 3790 1185
rect 3920 15 3940 1185
rect 4070 15 4090 1185
rect 4170 15 4190 1185
rect 4320 15 4340 1185
rect 4470 15 4490 1185
rect 4620 15 4640 1185
rect 4770 15 4790 1185
rect 4920 15 4940 1185
rect 5070 15 5090 1185
rect 5220 15 5240 1185
rect -190 -1495 -170 -325
rect -40 -1495 -20 -325
rect 110 -1495 130 -325
rect 190 -1495 210 -325
rect 340 -1495 360 -325
rect 490 -1495 510 -325
rect 640 -1495 660 -325
rect 790 -1495 810 -325
rect 940 -1495 960 -325
rect 1090 -1495 1110 -325
rect 1240 -1495 1260 -325
rect 1390 -1495 1410 -325
rect 1540 -1495 1560 -325
rect 1690 -1495 1710 -325
rect 1840 -1495 1860 -325
rect 1990 -1495 2010 -325
rect 2140 -1495 2160 -325
rect 2290 -1495 2310 -325
rect 2440 -1495 2460 -325
rect 2590 -1495 2610 -325
rect 2720 -1495 2740 -325
rect 2870 -1495 2890 -325
rect 2950 -1495 2970 -325
rect 3100 -1495 3120 -325
rect 3250 -1495 3270 -325
rect 3400 -1495 3420 -325
rect 3550 -1495 3570 -325
rect 3630 -1495 3650 -325
rect 3780 -1495 3800 -325
rect 3930 -1495 3950 -325
rect 4080 -1495 4100 -325
rect 4230 -1495 4250 -325
rect 4380 -1495 4400 -325
rect 4530 -1495 4550 -325
rect 4680 -1495 4700 -325
rect 4830 -1495 4850 -325
rect 4980 -1495 5000 -325
<< psubdiff >>
rect -255 1185 -205 1200
rect -255 15 -240 1185
rect -220 15 -205 1185
rect -255 0 -205 15
rect 1305 1185 1355 1200
rect 1305 15 1320 1185
rect 1340 15 1355 1185
rect 1305 0 1355 15
rect 4105 1185 4155 1200
rect 4105 15 4120 1185
rect 4140 15 4155 1185
rect 4105 0 4155 15
rect 5255 1185 5305 1200
rect 5255 15 5270 1185
rect 5290 15 5305 1185
rect 5255 0 5305 15
rect -255 -325 -205 -310
rect -255 -1495 -240 -325
rect -220 -1495 -205 -325
rect -255 -1510 -205 -1495
rect 2625 -325 2675 -310
rect 2625 -1495 2640 -325
rect 2660 -1495 2675 -325
rect 2625 -1510 2675 -1495
rect 5015 -325 5065 -310
rect 5015 -1495 5030 -325
rect 5050 -1495 5065 -325
rect 5015 -1510 5065 -1495
<< psubdiffcont >>
rect -240 15 -220 1185
rect 1320 15 1340 1185
rect 4120 15 4140 1185
rect 5270 15 5290 1185
rect -240 -1495 -220 -325
rect 2640 -1495 2660 -325
rect 5030 -1495 5050 -325
<< poly >>
rect 680 1240 720 1250
rect 680 1225 690 1240
rect 675 1220 690 1225
rect 710 1230 720 1240
rect 1705 1240 1745 1250
rect 1705 1230 1715 1240
rect 710 1220 1225 1230
rect 675 1215 1225 1220
rect 1555 1220 1715 1230
rect 1735 1230 1745 1240
rect 1915 1240 1955 1250
rect 1915 1230 1925 1240
rect 1735 1220 1925 1230
rect 1945 1230 1955 1240
rect 2560 1245 2600 1255
rect 2560 1235 2570 1245
rect 1945 1220 2405 1230
rect 1555 1215 2405 1220
rect -155 1200 -55 1215
rect -5 1200 95 1215
rect 145 1200 245 1215
rect 295 1200 395 1215
rect 445 1200 545 1215
rect 675 1200 775 1215
rect 825 1200 925 1215
rect 975 1200 1075 1215
rect 1125 1200 1225 1215
rect 1405 1200 1505 1215
rect 1555 1200 1655 1215
rect 1705 1200 1805 1215
rect 1855 1200 1955 1215
rect 2005 1200 2105 1215
rect 2155 1200 2255 1215
rect 2305 1200 2405 1215
rect 2455 1225 2570 1235
rect 2590 1235 2600 1245
rect 2860 1245 2900 1255
rect 2860 1235 2870 1245
rect 2590 1225 2870 1235
rect 2890 1235 2900 1245
rect 2990 1240 3370 1255
rect 2990 1235 3005 1240
rect 2890 1225 3005 1235
rect 2455 1215 3005 1225
rect 3355 1235 3370 1240
rect 3460 1245 3500 1255
rect 3460 1235 3470 1245
rect 3355 1225 3470 1235
rect 3490 1235 3500 1245
rect 3760 1245 3800 1255
rect 3760 1235 3770 1245
rect 3490 1225 3770 1235
rect 3790 1235 3800 1245
rect 4505 1240 4545 1250
rect 3790 1225 3905 1235
rect 4505 1230 4515 1240
rect 3355 1215 3905 1225
rect 2455 1200 2555 1215
rect 2605 1200 2705 1215
rect 2755 1200 2855 1215
rect 2905 1200 3005 1215
rect 3055 1200 3155 1215
rect 3205 1200 3305 1215
rect 3355 1200 3455 1215
rect 3505 1200 3605 1215
rect 3655 1200 3755 1215
rect 3805 1200 3905 1215
rect 3955 1220 4515 1230
rect 4535 1230 4545 1240
rect 4715 1240 4755 1250
rect 4715 1230 4725 1240
rect 4535 1220 4725 1230
rect 4745 1230 4755 1240
rect 4745 1220 4905 1230
rect 3955 1215 4905 1220
rect 3955 1200 4055 1215
rect 4205 1200 4305 1215
rect 4355 1200 4455 1215
rect 4505 1200 4605 1215
rect 4655 1200 4755 1215
rect 4805 1200 4905 1215
rect 4955 1200 5055 1215
rect 5105 1200 5205 1215
rect -155 -15 -55 0
rect -5 -10 95 0
rect 145 -10 245 0
rect 295 -10 395 0
rect 445 -10 545 0
rect -5 -20 545 -10
rect 675 -15 775 0
rect 825 -15 925 0
rect 975 -15 1075 0
rect 1125 -15 1225 0
rect 1405 -15 1505 0
rect 1555 -15 1655 0
rect 1705 -15 1805 0
rect 1855 -15 1955 0
rect 2005 -15 2105 0
rect 2155 -15 2255 0
rect 2305 -15 2405 0
rect 2455 -15 2555 0
rect 2605 -15 2705 0
rect 2755 -15 2855 0
rect 2905 -15 3005 0
rect 3055 -15 3155 0
rect -5 -25 260 -20
rect 250 -40 260 -25
rect 280 -25 545 -20
rect 1405 -20 1445 -15
rect 280 -40 290 -25
rect 250 -50 290 -40
rect 1405 -40 1415 -20
rect 1435 -40 1445 -20
rect 1405 -50 1445 -40
rect 2350 -20 2390 -15
rect 2350 -40 2360 -20
rect 2380 -40 2390 -20
rect 2350 -50 2390 -40
rect 250 -110 265 -50
rect 250 -120 290 -110
rect 250 -140 260 -120
rect 280 -140 290 -120
rect 250 -150 290 -140
rect 570 -140 610 -130
rect 570 -160 580 -140
rect 600 -155 610 -140
rect 690 -140 730 -130
rect 3140 -135 3155 -15
rect 690 -155 700 -140
rect 600 -160 700 -155
rect 720 -160 730 -140
rect 570 -170 730 -160
rect 3115 -145 3155 -135
rect 3115 -165 3125 -145
rect 3145 -165 3155 -145
rect 3115 -175 3155 -165
rect 3205 -15 3305 0
rect 3355 -15 3455 0
rect 3505 -15 3605 0
rect 3655 -15 3755 0
rect 3805 -15 3905 0
rect 3955 -15 4055 0
rect 4205 -15 4305 0
rect 4355 -15 4455 0
rect 4505 -15 4605 0
rect 4655 -15 4755 0
rect 4805 -15 4905 0
rect 4955 -15 5055 0
rect 5105 -15 5205 0
rect 3205 -135 3220 -15
rect 3205 -145 3245 -135
rect 3205 -165 3215 -145
rect 3235 -165 3245 -145
rect 3205 -175 3245 -165
rect 3655 -175 3670 -15
rect 3970 -20 4010 -15
rect 3970 -40 3980 -20
rect 4000 -40 4010 -20
rect 5015 -20 5055 -15
rect 5015 -40 5025 -20
rect 5045 -40 5055 -20
rect 3970 -50 4010 -40
rect 4400 -50 4560 -40
rect 5015 -50 5055 -40
rect 4400 -70 4410 -50
rect 4430 -55 4530 -50
rect 4430 -70 4440 -55
rect 4400 -80 4440 -70
rect 4520 -70 4530 -55
rect 4550 -70 4560 -50
rect 4520 -80 4560 -70
rect 4400 -115 4560 -105
rect 4400 -135 4410 -115
rect 4430 -120 4530 -115
rect 4430 -135 4440 -120
rect 4400 -145 4440 -135
rect 4520 -135 4530 -120
rect 4550 -135 4560 -115
rect 4520 -145 4560 -135
rect 3630 -185 3670 -175
rect 570 -205 730 -195
rect 570 -225 580 -205
rect 600 -210 700 -205
rect 600 -225 610 -210
rect 570 -235 610 -225
rect 690 -225 700 -210
rect 720 -225 730 -205
rect 3630 -205 3640 -185
rect 3660 -205 3670 -185
rect 3630 -215 3670 -205
rect 690 -235 730 -225
rect 330 -265 370 -255
rect 330 -280 340 -265
rect -5 -285 340 -280
rect 360 -280 370 -265
rect 630 -265 670 -255
rect 630 -280 640 -265
rect 360 -285 640 -280
rect 660 -280 670 -265
rect 930 -265 970 -255
rect 930 -280 940 -265
rect 660 -285 940 -280
rect 960 -280 970 -265
rect 1230 -265 1270 -255
rect 1230 -280 1240 -265
rect 960 -285 1240 -280
rect 1260 -280 1270 -265
rect 1530 -265 1570 -255
rect 1530 -280 1540 -265
rect 1260 -285 1540 -280
rect 1560 -280 1570 -265
rect 1830 -265 1870 -255
rect 1830 -280 1840 -265
rect 1560 -285 1840 -280
rect 1860 -280 1870 -265
rect 2130 -265 2170 -255
rect 2130 -280 2140 -265
rect 1860 -285 2140 -280
rect 2160 -280 2170 -265
rect 2430 -265 2470 -255
rect 2430 -280 2440 -265
rect 2160 -285 2440 -280
rect 2460 -280 2470 -265
rect 3090 -265 3130 -255
rect 3090 -280 3100 -265
rect 2460 -285 2855 -280
rect -5 -295 2855 -285
rect -155 -310 -55 -295
rect -5 -310 95 -295
rect 225 -310 325 -295
rect 375 -310 475 -295
rect 525 -310 625 -295
rect 675 -310 775 -295
rect 825 -310 925 -295
rect 975 -310 1075 -295
rect 1125 -310 1225 -295
rect 1275 -310 1375 -295
rect 1425 -310 1525 -295
rect 1575 -310 1675 -295
rect 1725 -310 1825 -295
rect 1875 -310 1975 -295
rect 2025 -310 2125 -295
rect 2175 -310 2275 -295
rect 2325 -310 2425 -295
rect 2475 -310 2575 -295
rect 2755 -310 2855 -295
rect 2985 -285 3100 -280
rect 3120 -280 3130 -265
rect 3390 -265 3430 -255
rect 3390 -280 3400 -265
rect 3120 -285 3400 -280
rect 3420 -280 3430 -265
rect 3680 -265 3720 -255
rect 3680 -280 3690 -265
rect 3420 -285 3535 -280
rect 2985 -295 3535 -285
rect 2985 -310 3085 -295
rect 3135 -310 3235 -295
rect 3285 -310 3385 -295
rect 3435 -310 3535 -295
rect 3665 -285 3690 -280
rect 3710 -280 3720 -265
rect 3710 -285 4815 -280
rect 3665 -295 4815 -285
rect 3665 -310 3765 -295
rect 3815 -310 3915 -295
rect 3965 -310 4065 -295
rect 4115 -310 4215 -295
rect 4265 -310 4365 -295
rect 4415 -310 4515 -295
rect 4565 -310 4665 -295
rect 4715 -310 4815 -295
rect 4865 -310 4965 -295
rect -155 -1525 -55 -1510
rect -5 -1525 95 -1510
rect 225 -1525 325 -1510
rect 375 -1525 475 -1510
rect 525 -1525 625 -1510
rect 675 -1525 775 -1510
rect 825 -1525 925 -1510
rect 975 -1525 1075 -1510
rect 1125 -1525 1225 -1510
rect 1275 -1525 1375 -1510
rect 1425 -1525 1525 -1510
rect 1575 -1525 1675 -1510
rect 1725 -1525 1825 -1510
rect 1875 -1525 1975 -1510
rect 2025 -1525 2125 -1510
rect 2175 -1525 2275 -1510
rect 2325 -1525 2425 -1510
rect 2475 -1525 2575 -1510
rect 2755 -1525 2855 -1510
rect 2985 -1525 3085 -1510
rect 3135 -1525 3235 -1510
rect 3285 -1525 3385 -1510
rect 3435 -1525 3535 -1510
rect 3665 -1525 3765 -1510
rect 3815 -1525 3915 -1510
rect 3965 -1525 4065 -1510
rect 4115 -1525 4215 -1510
rect 4265 -1525 4365 -1510
rect 4415 -1525 4515 -1510
rect 4565 -1525 4665 -1510
rect 4715 -1525 4815 -1510
rect 4865 -1525 4965 -1510
<< polycont >>
rect 690 1220 710 1240
rect 1715 1220 1735 1240
rect 1925 1220 1945 1240
rect 2570 1225 2590 1245
rect 2870 1225 2890 1245
rect 3470 1225 3490 1245
rect 3770 1225 3790 1245
rect 4515 1220 4535 1240
rect 4725 1220 4745 1240
rect 260 -40 280 -20
rect 1415 -40 1435 -20
rect 2360 -40 2380 -20
rect 260 -140 280 -120
rect 580 -160 600 -140
rect 700 -160 720 -140
rect 3125 -165 3145 -145
rect 3215 -165 3235 -145
rect 3980 -40 4000 -20
rect 5025 -40 5045 -20
rect 4410 -70 4430 -50
rect 4530 -70 4550 -50
rect 4410 -135 4430 -115
rect 4530 -135 4550 -115
rect 580 -225 600 -205
rect 700 -225 720 -205
rect 3640 -205 3660 -185
rect 340 -285 360 -265
rect 640 -285 660 -265
rect 940 -285 960 -265
rect 1240 -285 1260 -265
rect 1540 -285 1560 -265
rect 1840 -285 1860 -265
rect 2140 -285 2160 -265
rect 2440 -285 2460 -265
rect 3100 -285 3120 -265
rect 3400 -285 3420 -265
rect 3690 -285 3710 -265
<< locali >>
rect 680 1240 720 1250
rect 550 1220 690 1240
rect 710 1220 720 1240
rect 550 1215 720 1220
rect -250 1185 -160 1195
rect -250 15 -240 1185
rect -220 15 -190 1185
rect -170 15 -160 1185
rect -250 5 -160 15
rect -50 1185 -10 1195
rect -50 15 -40 1185
rect -20 15 -10 1185
rect -50 -70 -10 15
rect 100 1185 140 1195
rect 100 15 110 1185
rect 130 15 140 1185
rect 100 5 140 15
rect 250 1185 290 1195
rect 250 15 260 1185
rect 280 15 290 1185
rect 250 -20 290 15
rect 400 1185 440 1195
rect 400 15 410 1185
rect 430 15 440 1185
rect 400 5 440 15
rect 550 1185 590 1215
rect 680 1210 720 1215
rect 1660 1240 1745 1250
rect 1660 1220 1715 1240
rect 1735 1220 1745 1240
rect 1660 1210 1745 1220
rect 1915 1240 2000 1250
rect 1915 1220 1925 1240
rect 1945 1220 2000 1240
rect 1915 1210 2000 1220
rect 550 15 560 1185
rect 580 15 590 1185
rect 250 -40 260 -20
rect 280 -40 290 -20
rect 250 -50 290 -40
rect 550 -70 590 15
rect -50 -90 590 -70
rect 250 -120 290 -110
rect 250 -140 260 -120
rect 280 -140 290 -120
rect 250 -150 290 -140
rect 570 -130 590 -90
rect 630 1185 670 1195
rect 630 15 640 1185
rect 660 15 670 1185
rect 630 -40 670 15
rect 780 1185 820 1195
rect 780 15 790 1185
rect 810 15 820 1185
rect 780 5 820 15
rect 930 1185 970 1195
rect 930 15 940 1185
rect 960 15 970 1185
rect 930 5 970 15
rect 1080 1185 1120 1195
rect 1080 15 1090 1185
rect 1110 15 1120 1185
rect 1080 5 1120 15
rect 1230 1185 1270 1195
rect 1230 15 1240 1185
rect 1260 15 1270 1185
rect 1230 -40 1270 15
rect 1310 1185 1400 1195
rect 1310 15 1320 1185
rect 1340 15 1370 1185
rect 1390 15 1400 1185
rect 1310 5 1400 15
rect 630 -60 1270 -40
rect 1360 -10 1400 5
rect 1510 1185 1550 1195
rect 1510 15 1520 1185
rect 1540 15 1550 1185
rect 1360 -20 1445 -10
rect 1360 -40 1415 -20
rect 1435 -40 1445 -20
rect 1360 -50 1445 -40
rect 570 -140 610 -130
rect 250 -215 270 -150
rect 570 -160 580 -140
rect 600 -160 610 -140
rect 570 -170 610 -160
rect 570 -205 610 -195
rect 570 -215 580 -205
rect -50 -225 580 -215
rect 600 -225 610 -205
rect -50 -235 610 -225
rect -50 -315 -10 -235
rect 330 -265 370 -255
rect 330 -285 340 -265
rect 360 -285 370 -265
rect -250 -325 -160 -315
rect -250 -1495 -240 -325
rect -220 -1495 -190 -325
rect -170 -1495 -160 -325
rect -250 -1505 -160 -1495
rect -55 -325 -10 -315
rect -55 -1495 -40 -325
rect -20 -1495 -10 -325
rect -55 -1505 -10 -1495
rect 100 -325 140 -315
rect 100 -1495 110 -325
rect 130 -1495 140 -325
rect 100 -1500 140 -1495
rect 180 -325 220 -315
rect 180 -1495 190 -325
rect 210 -1495 220 -325
rect 180 -1525 220 -1495
rect 330 -325 370 -285
rect 630 -265 670 -60
rect 1425 -95 1445 -50
rect 1510 -55 1550 15
rect 1660 1185 1700 1210
rect 1660 15 1670 1185
rect 1690 15 1700 1185
rect 1660 5 1700 15
rect 1810 1185 1850 1195
rect 1810 15 1820 1185
rect 1840 15 1850 1185
rect 1810 -55 1850 15
rect 1960 1185 2000 1210
rect 2560 1245 2600 1255
rect 2560 1225 2570 1245
rect 2590 1225 2600 1245
rect 1960 15 1970 1185
rect 1990 15 2000 1185
rect 1960 5 2000 15
rect 2110 1185 2150 1195
rect 2110 15 2120 1185
rect 2140 15 2150 1185
rect 2110 -55 2150 15
rect 2260 1185 2300 1195
rect 2260 15 2270 1185
rect 2290 15 2300 1185
rect 2260 5 2300 15
rect 2410 1185 2450 1195
rect 2410 15 2420 1185
rect 2440 15 2450 1185
rect 2350 -20 2390 -10
rect 2350 -40 2360 -20
rect 2380 -40 2390 -20
rect 2410 -15 2450 15
rect 2560 1185 2600 1225
rect 2860 1245 2900 1255
rect 2860 1225 2870 1245
rect 2890 1225 2900 1245
rect 2560 15 2570 1185
rect 2590 15 2600 1185
rect 2560 5 2600 15
rect 2710 1185 2750 1195
rect 2710 15 2720 1185
rect 2740 15 2750 1185
rect 2710 -15 2750 15
rect 2860 1185 2900 1225
rect 3460 1245 3500 1255
rect 3460 1225 3470 1245
rect 3490 1225 3500 1245
rect 2860 15 2870 1185
rect 2890 15 2900 1185
rect 2860 5 2900 15
rect 3010 1185 3050 1195
rect 3010 15 3020 1185
rect 3040 15 3050 1185
rect 3010 -15 3050 15
rect 3160 1185 3200 1195
rect 3160 15 3170 1185
rect 3190 15 3200 1185
rect 3160 5 3200 15
rect 3310 1185 3350 1195
rect 3310 15 3320 1185
rect 3340 15 3350 1185
rect 3310 -15 3350 15
rect 3460 1185 3500 1225
rect 3760 1245 3800 1255
rect 3760 1225 3770 1245
rect 3790 1225 3800 1245
rect 3460 15 3470 1185
rect 3490 15 3500 1185
rect 3460 5 3500 15
rect 3610 1185 3650 1195
rect 3610 15 3620 1185
rect 3640 15 3650 1185
rect 3610 -15 3650 15
rect 3760 1185 3800 1225
rect 4460 1240 4545 1250
rect 4460 1220 4515 1240
rect 4535 1220 4545 1240
rect 4460 1210 4545 1220
rect 4715 1240 4800 1250
rect 4715 1220 4725 1240
rect 4745 1220 4800 1240
rect 4715 1210 4800 1220
rect 3760 15 3770 1185
rect 3790 15 3800 1185
rect 3760 5 3800 15
rect 3910 1185 3950 1195
rect 3910 15 3920 1185
rect 3940 15 3950 1185
rect 3910 -15 3950 15
rect 4060 1185 4200 1195
rect 4060 15 4070 1185
rect 4090 15 4120 1185
rect 4140 15 4170 1185
rect 4190 15 4200 1185
rect 4060 5 4200 15
rect 4310 1185 4350 1195
rect 4310 15 4320 1185
rect 4340 15 4350 1185
rect 2410 -35 3950 -15
rect 3970 -20 4010 -10
rect 2350 -50 2390 -40
rect 2370 -55 2390 -50
rect 3970 -40 3980 -20
rect 4000 -40 4010 -20
rect 3970 -50 4010 -40
rect 3970 -55 3990 -50
rect 4310 -55 4350 15
rect 4460 1185 4500 1210
rect 4460 15 4470 1185
rect 4490 15 4500 1185
rect 4400 -50 4440 -40
rect 4400 -55 4410 -50
rect 1510 -75 2330 -55
rect 2370 -75 3990 -55
rect 4030 -70 4410 -55
rect 4430 -70 4440 -50
rect 4030 -75 4440 -70
rect 2310 -95 2330 -75
rect 4030 -95 4050 -75
rect 4400 -80 4440 -75
rect 1425 -115 2290 -95
rect 2310 -115 4050 -95
rect 4070 -115 4440 -105
rect 690 -140 730 -130
rect 690 -160 700 -140
rect 720 -150 730 -140
rect 2270 -135 2290 -115
rect 4070 -125 4410 -115
rect 4070 -135 4090 -125
rect 2270 -145 4090 -135
rect 4400 -135 4410 -125
rect 4430 -135 4440 -115
rect 4400 -145 4440 -135
rect 720 -160 770 -150
rect 2270 -155 3125 -145
rect 690 -170 770 -160
rect 750 -175 770 -170
rect 3115 -165 3125 -155
rect 3145 -155 3215 -145
rect 3145 -165 3155 -155
rect 3115 -175 3155 -165
rect 3205 -165 3215 -155
rect 3235 -155 4090 -145
rect 3235 -165 3245 -155
rect 3205 -175 3245 -165
rect 750 -195 2980 -175
rect 690 -205 730 -195
rect 690 -225 700 -205
rect 720 -215 730 -205
rect 2940 -215 2980 -195
rect 3620 -185 3670 -175
rect 3620 -205 3640 -185
rect 3660 -205 3670 -185
rect 3620 -215 3670 -205
rect 720 -225 2900 -215
rect 690 -235 2900 -225
rect 630 -285 640 -265
rect 660 -285 670 -265
rect 330 -1495 340 -325
rect 360 -1495 370 -325
rect 330 -1505 370 -1495
rect 480 -325 520 -315
rect 480 -1495 490 -325
rect 510 -1495 520 -325
rect 480 -1525 520 -1495
rect 630 -325 670 -285
rect 930 -265 970 -255
rect 930 -285 940 -265
rect 960 -285 970 -265
rect 630 -1495 640 -325
rect 660 -1495 670 -325
rect 630 -1505 670 -1495
rect 780 -325 820 -315
rect 780 -1495 790 -325
rect 810 -1495 820 -325
rect 780 -1525 820 -1495
rect 930 -325 970 -285
rect 1230 -265 1270 -255
rect 1230 -285 1240 -265
rect 1260 -285 1270 -265
rect 930 -1495 940 -325
rect 960 -1495 970 -325
rect 930 -1505 970 -1495
rect 1080 -325 1120 -315
rect 1080 -1495 1090 -325
rect 1110 -1495 1120 -325
rect 1080 -1525 1120 -1495
rect 1230 -325 1270 -285
rect 1530 -265 1570 -255
rect 1530 -285 1540 -265
rect 1560 -285 1570 -265
rect 1230 -1495 1240 -325
rect 1260 -1495 1270 -325
rect 1230 -1505 1270 -1495
rect 1380 -325 1420 -315
rect 1380 -1495 1390 -325
rect 1410 -1495 1420 -325
rect 1380 -1525 1420 -1495
rect 1530 -325 1570 -285
rect 1830 -265 1870 -255
rect 1830 -285 1840 -265
rect 1860 -285 1870 -265
rect 1530 -1495 1540 -325
rect 1560 -1495 1570 -325
rect 1530 -1505 1570 -1495
rect 1680 -325 1720 -315
rect 1680 -1495 1690 -325
rect 1710 -1495 1720 -325
rect 1680 -1525 1720 -1495
rect 1830 -325 1870 -285
rect 2130 -265 2170 -255
rect 2130 -285 2140 -265
rect 2160 -285 2170 -265
rect 1830 -1495 1840 -325
rect 1860 -1495 1870 -325
rect 1830 -1505 1870 -1495
rect 1980 -325 2020 -315
rect 1980 -1495 1990 -325
rect 2010 -1495 2020 -325
rect 1980 -1525 2020 -1495
rect 2130 -325 2170 -285
rect 2430 -265 2470 -255
rect 2430 -285 2440 -265
rect 2460 -285 2470 -265
rect 2130 -1495 2140 -325
rect 2160 -1495 2170 -325
rect 2130 -1505 2170 -1495
rect 2280 -325 2320 -315
rect 2280 -1495 2290 -325
rect 2310 -1495 2320 -325
rect 2280 -1525 2320 -1495
rect 2430 -325 2470 -285
rect 2430 -1495 2440 -325
rect 2460 -1495 2470 -325
rect 2430 -1505 2470 -1495
rect 2580 -325 2670 -315
rect 2580 -1495 2590 -325
rect 2610 -1495 2640 -325
rect 2660 -1495 2670 -325
rect 2580 -1505 2670 -1495
rect 2710 -325 2750 -315
rect 2710 -1495 2720 -325
rect 2740 -1495 2750 -325
rect 2710 -1505 2750 -1495
rect 2860 -325 2900 -235
rect 2860 -1495 2870 -325
rect 2890 -1495 2900 -325
rect 2860 -1505 2900 -1495
rect 2940 -235 3580 -215
rect 2940 -325 2980 -235
rect 2940 -1495 2950 -325
rect 2970 -1495 2980 -325
rect 2940 -1505 2980 -1495
rect 3090 -265 3130 -255
rect 3090 -285 3100 -265
rect 3120 -285 3130 -265
rect 3090 -325 3130 -285
rect 3390 -265 3430 -255
rect 3390 -285 3400 -265
rect 3420 -285 3430 -265
rect 3090 -1495 3100 -325
rect 3120 -1495 3130 -325
rect 3090 -1505 3130 -1495
rect 3240 -325 3280 -315
rect 3240 -1495 3250 -325
rect 3270 -1495 3280 -325
rect 3240 -1505 3280 -1495
rect 3390 -325 3430 -285
rect 3390 -1495 3400 -325
rect 3420 -1495 3430 -325
rect 3390 -1505 3430 -1495
rect 3540 -325 3580 -235
rect 3540 -1495 3550 -325
rect 3570 -1495 3580 -325
rect 3540 -1505 3580 -1495
rect 3620 -325 3660 -215
rect 3680 -265 3720 -255
rect 4460 -260 4500 15
rect 4610 1185 4650 1195
rect 4610 15 4620 1185
rect 4640 15 4650 1185
rect 4520 -50 4560 -40
rect 4520 -70 4530 -50
rect 4550 -55 4560 -50
rect 4610 -55 4650 15
rect 4760 1185 4800 1210
rect 4760 15 4770 1185
rect 4790 15 4800 1185
rect 4760 5 4800 15
rect 4910 1185 4950 1195
rect 4910 15 4920 1185
rect 4940 15 4950 1185
rect 4910 -55 4950 15
rect 5060 1185 5100 1195
rect 5060 15 5070 1185
rect 5090 15 5100 1185
rect 5060 -10 5100 15
rect 5210 1185 5300 1195
rect 5210 15 5220 1185
rect 5240 15 5270 1185
rect 5290 15 5300 1185
rect 5210 5 5300 15
rect 4550 -70 4950 -55
rect 4520 -75 4950 -70
rect 5015 -20 5100 -10
rect 5015 -40 5025 -20
rect 5045 -40 5100 -20
rect 5015 -50 5100 -40
rect 4520 -80 4560 -75
rect 5015 -105 5035 -50
rect 4520 -115 5035 -105
rect 4520 -135 4530 -115
rect 4550 -125 5035 -115
rect 4550 -135 4560 -125
rect 4520 -145 4560 -135
rect 3680 -285 3690 -265
rect 3710 -285 3720 -265
rect 3680 -295 3720 -285
rect 4220 -280 4500 -260
rect 3620 -1495 3630 -325
rect 3650 -1495 3660 -325
rect 2580 -1525 2620 -1505
rect 180 -1545 2620 -1525
rect 3620 -1525 3660 -1495
rect 3770 -325 3810 -315
rect 3770 -1495 3780 -325
rect 3800 -1495 3810 -325
rect 3770 -1505 3810 -1495
rect 3920 -325 3960 -315
rect 3920 -1495 3930 -325
rect 3950 -1495 3960 -325
rect 3920 -1505 3960 -1495
rect 4070 -325 4110 -315
rect 4070 -1495 4080 -325
rect 4100 -1495 4110 -325
rect 4070 -1505 4110 -1495
rect 4220 -325 4260 -280
rect 4220 -1495 4230 -325
rect 4250 -1495 4260 -325
rect 4220 -1505 4260 -1495
rect 4370 -325 4410 -315
rect 4370 -1495 4380 -325
rect 4400 -1495 4410 -325
rect 4370 -1505 4410 -1495
rect 4520 -325 4560 -315
rect 4520 -1495 4530 -325
rect 4550 -1495 4560 -325
rect 4520 -1505 4560 -1495
rect 4670 -325 4710 -315
rect 4670 -1495 4680 -325
rect 4700 -1495 4710 -325
rect 4670 -1505 4710 -1495
rect 4820 -325 4860 -315
rect 4820 -1495 4830 -325
rect 4850 -1495 4860 -325
rect 4820 -1525 4860 -1495
rect 4970 -325 5060 -315
rect 4970 -1495 4980 -325
rect 5000 -1495 5030 -325
rect 5050 -1495 5060 -325
rect 4970 -1505 5060 -1495
rect 3620 -1545 4860 -1525
<< viali >>
rect 790 15 810 1185
rect 940 15 960 1185
rect 3100 -285 3120 -265
<< metal1 >>
rect 780 1190 820 1195
rect 780 10 785 1190
rect 815 10 820 1190
rect 780 5 820 10
rect 930 1185 970 1195
rect 930 15 940 1185
rect 960 15 970 1185
rect 930 -135 970 15
rect 930 -175 5335 -135
rect 3090 -265 3130 -175
rect 3090 -285 3100 -265
rect 3120 -285 3130 -265
rect 3090 -295 3130 -285
<< via1 >>
rect 785 1185 815 1190
rect 785 15 790 1185
rect 790 15 810 1185
rect 810 15 815 1185
rect 785 10 815 15
<< metal2 >>
rect 780 1190 820 1195
rect 780 10 785 1190
rect 815 10 820 1190
rect 780 5 820 10
<< end >>
