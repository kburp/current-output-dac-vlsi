* NGSPICE file created from big.ext - technology: sky130A


* Top level circuit big

X0 a_9330_n3020# VBN VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X1 a_n10_n3050# a_n10_n3050# ROUT VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X2 VBN VBN VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X3 a_n110_0# VP VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=1
X4 a_n110_n3020# VN VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=1
X5 ROUT a_n10_n3050# a_n10_n3050# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X6 VBN a_n110_0# VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X7 a_n10_n3050# a_n110_0# VP VP sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=1
X8 a_n10_n3050# a_n10_n3050# ROUT VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X9 a_2910_0# VIN VIN VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=1
X10 a_5010_n30# a_5010_n30# a_4910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X11 a_n110_n3020# a_n10_n3050# VN VN sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=6 ps=25 w=12 l=1
X12 a_2910_0# a_3010_n30# a_3010_n30# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X13 ROUT a_n10_n3050# a_n10_n3050# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X14 a_n10_n3050# a_n10_n3050# ROUT VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X15 a_5010_n30# a_5010_n30# a_4910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X16 VOUT VIN a_4910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X17 ROUT a_n10_n3050# a_n10_n3050# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X18 a_2910_0# a_3010_n30# a_3010_n30# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X19 a_2910_0# a_3010_n30# VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=1
X20 a_8130_n3020# VBN VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X21 VP a_n110_n3020# a_n110_n3020# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X22 a_5010_n30# a_5010_n30# a_4910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X23 a_2910_0# a_3010_n30# a_3010_n30# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X24 VP VP VIN VP sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=1
X25 a_n10_n3050# a_n10_n3050# ROUT VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X26 a_5010_n30# a_5010_n30# a_4910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X27 VN VBN a_n110_0# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=1
X28 VN VBN a_8730_n3020# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X29 VP a_3010_n30# a_4910_0# VP sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=1
X30 a_2910_0# a_3010_n30# a_3010_n30# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X31 ROUT a_n10_n3050# a_n10_n3050# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X32 a_n110_0# VBN VN VN sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=1
X33 VN VN a_5010_n30# VN sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=1
X34 VN a_n10_n3050# a_n110_n3020# VN sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=1
X35 a_n10_n3050# a_n10_n3050# ROUT VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=1
X36 ROUT a_n10_n3050# a_n10_n3050# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X37 VP a_n110_n3020# a_n110_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X38 a_n10_n3050# a_n10_n3050# ROUT VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X39 VN VBN a_7530_n3020# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X40 VP a_n110_0# a_n10_n3050# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=1
X41 ROUT a_n10_n3050# a_n10_n3050# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X42 a_8730_n3020# VBN a_3010_n30# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X43 VP a_n110_0# VBN VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X44 a_3010_n30# a_3010_n30# a_2910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X45 a_4910_0# a_3010_n30# VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=1
X46 a_n10_n3050# a_n10_n3050# ROUT VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X47 a_4910_0# a_5010_n30# a_5010_n30# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X48 VN VBN VBN VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X49 a_5010_n30# VBN a_9330_n3020# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X50 a_3010_n30# a_3010_n30# a_2910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X51 a_n10_n3050# a_n10_n3050# ROUT VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X52 VP a_3010_n30# a_2910_0# VP sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=1
X53 a_4910_0# a_5010_n30# a_5010_n30# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X54 a_n110_n3020# a_n110_n3020# VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X55 a_4910_0# VIN VOUT VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X56 VIN VIN a_2910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X57 a_4910_0# a_5010_n30# a_5010_n30# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X58 a_3010_n30# a_3010_n30# a_2910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X59 a_7530_n3020# VBN a_5010_n30# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=1
X60 a_n110_0# a_n110_n3020# VP VP sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=1
X61 a_3010_n30# a_3010_n30# a_2910_0# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X62 ROUT a_n10_n3050# a_n10_n3050# VN sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=1
X63 a_4910_0# a_5010_n30# a_5010_n30# VP sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X64 a_3010_n30# VBN a_8130_n3020# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
X65 ROUT a_n10_n3050# a_n10_n3050# VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=1
.end

