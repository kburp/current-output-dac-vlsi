* NGSPICE file created from dac.ext - technology: sky130A


* Top level circuit dac

X0 a_3500_n4800# Vgate a_2300_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X1 a_3500_n4800# b3 VN VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X2 a_200_400# Vgate a_1100_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X3 Iout Vgate a_200_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X4 a_200_n4800# Vgate a_1100_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X5 a_2300_400# Vgate a_500_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X6 VN b0 a_200_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X7 a_2300_400# Vgate a_1100_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X8 a_2300_n4800# Vgate a_1100_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X9 a_200_400# VN VN VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=12 ps=49 w=24 l=1
X10 a_500_400# Vgate a_2300_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X11 a_2300_n4800# Vgate a_1100_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X12 a_500_400# b1 VN VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X13 a_3500_n4800# Vgate a_2300_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X14 a_1100_400# Vgate a_500_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X15 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=96 ps=392 w=24 l=1
X16 a_2300_400# Vgate a_3500_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X17 a_200_n4800# VN VN VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=12 ps=49 w=24 l=1
X18 VN b4 a_2300_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X19 VN b2 a_2300_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X20 VN VN a_1100_400# VN sky130_fd_pr__nfet_01v8 ad=12 pd=49 as=6 ps=24.5 w=24 l=1
X21 VP a_1100_400# a_1100_400# VP sky130_fd_pr__pfet_01v8 ad=12 pd=49 as=12 ps=49 w=24 l=1
X22 a_1100_n4800# b5 VN VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X23 a_1100_n4800# Vgate a_200_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X24 a_1100_400# Vgate a_1100_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X25 a_500_400# Vgate a_200_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X26 a_2300_n4800# Vgate a_3500_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X27 a_1100_400# Vgate a_3500_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X28 a_200_400# Vgate a_500_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X29 a_200_n4800# Vgate Iout VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X30 VN b6 a_200_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X31 a_1100_400# Vgate a_200_400# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
X32 a_1100_n4800# Vgate a_2300_n4800# VN sky130_fd_pr__nfet_01v8 ad=6 pd=24.5 as=6 ps=24.5 w=24 l=1
.end

