magic
tech sky130A
timestamp 1699649434
<< nwell >>
rect 75 120 295 395
<< nmos >>
rect 145 -15 160 85
rect 210 -15 225 85
rect 210 -150 225 -50
<< pmos >>
rect 210 275 225 375
rect 145 140 160 240
rect 210 140 225 240
<< ndiff >>
rect 95 70 145 85
rect 95 0 110 70
rect 130 0 145 70
rect 95 -15 145 0
rect 160 70 210 85
rect 160 0 175 70
rect 195 0 210 70
rect 160 -15 210 0
rect 225 70 275 85
rect 225 0 240 70
rect 260 0 275 70
rect 225 -15 275 0
rect 160 -65 210 -50
rect 160 -135 175 -65
rect 195 -135 210 -65
rect 160 -150 210 -135
rect 225 -65 275 -50
rect 225 -135 240 -65
rect 260 -135 275 -65
rect 225 -150 275 -135
<< pdiff >>
rect 160 360 210 375
rect 160 290 175 360
rect 195 290 210 360
rect 160 275 210 290
rect 225 360 275 375
rect 225 290 240 360
rect 260 290 275 360
rect 225 275 275 290
rect 95 225 145 240
rect 95 155 110 225
rect 130 155 145 225
rect 95 140 145 155
rect 160 225 210 240
rect 160 155 175 225
rect 195 155 210 225
rect 160 140 210 155
rect 225 225 275 240
rect 225 155 240 225
rect 260 155 275 225
rect 225 140 275 155
<< ndiffc >>
rect 110 0 130 70
rect 175 0 195 70
rect 240 0 260 70
rect 175 -135 195 -65
rect 240 -135 260 -65
<< pdiffc >>
rect 175 290 195 360
rect 240 290 260 360
rect 110 155 130 225
rect 175 155 195 225
rect 240 155 260 225
<< poly >>
rect 210 375 225 390
rect 105 310 145 320
rect 105 290 115 310
rect 135 290 145 310
rect 105 280 145 290
rect 130 265 145 280
rect 130 250 160 265
rect 145 240 160 250
rect 210 240 225 275
rect 145 85 160 140
rect 210 85 225 140
rect 145 -25 160 -15
rect 130 -40 160 -25
rect 130 -55 145 -40
rect 210 -50 225 -15
rect 105 -65 145 -55
rect 105 -85 115 -65
rect 135 -85 145 -65
rect 105 -95 145 -85
rect 210 -165 225 -150
<< polycont >>
rect 115 290 135 310
rect 115 -85 135 -65
<< locali >>
rect 165 360 205 370
rect 165 320 175 360
rect 105 310 175 320
rect 105 290 115 310
rect 135 290 175 310
rect 195 290 205 360
rect 105 280 205 290
rect 230 360 270 370
rect 230 290 240 360
rect 260 290 270 360
rect 230 280 270 290
rect 100 225 140 235
rect 100 155 110 225
rect 130 155 140 225
rect 100 145 140 155
rect 165 225 205 235
rect 165 155 175 225
rect 195 155 205 225
rect 100 70 140 80
rect 100 0 110 70
rect 130 0 140 70
rect 100 -10 140 0
rect 165 70 205 155
rect 230 225 270 235
rect 230 155 240 225
rect 260 155 270 225
rect 230 145 270 155
rect 165 0 175 70
rect 195 0 205 70
rect 165 -10 205 0
rect 230 70 270 80
rect 230 0 240 70
rect 260 0 270 70
rect 230 -10 270 0
rect 105 -65 205 -55
rect 105 -85 115 -65
rect 135 -85 175 -65
rect 105 -95 175 -85
rect 165 -135 175 -95
rect 195 -135 205 -65
rect 165 -145 205 -135
rect 230 -65 270 -55
rect 230 -135 240 -65
rect 260 -135 270 -65
rect 230 -145 270 -135
<< viali >>
rect 240 290 260 360
rect 110 155 130 225
rect 110 0 130 70
rect 240 155 260 225
rect 240 0 260 70
rect 240 -135 260 -65
<< metal1 >>
rect 230 365 270 370
rect 230 285 235 365
rect 265 285 270 365
rect 230 280 270 285
rect 100 225 140 235
rect 100 155 110 225
rect 130 155 140 225
rect 100 145 140 155
rect 230 230 270 235
rect 230 150 235 230
rect 265 150 270 230
rect 230 145 270 150
rect 120 120 140 145
rect 120 100 250 120
rect 230 80 250 100
rect 100 75 140 80
rect 100 -5 105 75
rect 135 -5 140 75
rect 100 -10 140 -5
rect 230 70 270 80
rect 230 0 240 70
rect 260 0 270 70
rect 230 -10 270 0
rect 230 -60 270 -55
rect 230 -140 235 -60
rect 265 -140 270 -60
rect 230 -145 270 -140
<< via1 >>
rect 235 360 265 365
rect 235 290 240 360
rect 240 290 260 360
rect 260 290 265 360
rect 235 285 265 290
rect 235 225 265 230
rect 235 155 240 225
rect 240 155 260 225
rect 260 155 265 225
rect 235 150 265 155
rect 105 70 135 75
rect 105 0 110 70
rect 110 0 130 70
rect 130 0 135 70
rect 105 -5 135 0
rect 235 -65 265 -60
rect 235 -135 240 -65
rect 240 -135 260 -65
rect 260 -135 265 -65
rect 235 -140 265 -135
<< metal2 >>
rect 230 365 270 370
rect 230 285 235 365
rect 265 285 270 365
rect 230 280 270 285
rect 230 230 270 235
rect 230 150 235 230
rect 265 150 270 230
rect 230 80 270 150
rect 100 75 270 80
rect 100 -5 105 75
rect 135 -5 270 75
rect 100 -10 270 -5
rect 230 -60 270 -10
rect 230 -140 235 -60
rect 265 -140 270 -60
rect 230 -145 270 -140
<< labels >>
rlabel metal2 270 100 270 100 3 VN
port 2 e
rlabel metal1 120 110 120 110 7 Vbn
port 3 w
rlabel metal2 270 325 270 325 3 VP
port 4 e
rlabel locali 205 95 205 95 3 Y
port 1 e
<< end >>
