magic
tech sky130A
timestamp 1699554853
<< nmos >>
rect 0 0 100 2400
rect 150 0 250 2400
rect 300 0 400 2400
rect 450 0 550 2400
rect 600 0 700 2400
rect 750 0 850 2400
rect 900 0 1000 2400
rect 1050 0 1150 2400
rect 1200 0 1300 2400
rect 1350 0 1450 2400
rect 1500 0 1600 2400
rect 1650 0 1750 2400
rect 1800 0 1900 2400
rect 1950 0 2050 2400
rect 2100 0 2200 2400
rect 2250 0 2350 2400
<< ndiff >>
rect -50 2385 0 2400
rect -50 15 -40 2385
rect -15 15 0 2385
rect -50 0 0 15
rect 100 0 150 2400
rect 250 0 300 2400
rect 400 0 450 2400
rect 550 0 600 2400
rect 700 0 750 2400
rect 850 0 900 2400
rect 1000 0 1050 2400
rect 1150 0 1200 2400
rect 1300 0 1350 2400
rect 1450 0 1500 2400
rect 1600 0 1650 2400
rect 1750 0 1800 2400
rect 1900 0 1950 2400
rect 2050 0 2100 2400
rect 2200 0 2250 2400
rect 2350 2385 2400 2400
rect 2350 15 2365 2385
rect 2390 15 2400 2385
rect 2350 0 2400 15
<< ndiffc >>
rect -40 15 -15 2385
rect 2365 15 2390 2385
<< psubdiff >>
rect -100 2385 -50 2400
rect -100 15 -85 2385
rect -60 15 -50 2385
rect -100 0 -50 15
rect 2400 2385 2450 2400
rect 2400 15 2410 2385
rect 2435 15 2450 2385
rect 2400 0 2450 15
<< psubdiffcont >>
rect -85 15 -60 2385
rect 2410 15 2435 2385
<< poly >>
rect 0 2400 100 2415
rect 150 2400 250 2415
rect 300 2400 400 2415
rect 450 2400 550 2415
rect 600 2400 700 2415
rect 750 2400 850 2415
rect 900 2400 1000 2415
rect 1050 2400 1150 2415
rect 1200 2400 1300 2415
rect 1350 2400 1450 2415
rect 1500 2400 1600 2415
rect 1650 2400 1750 2415
rect 1800 2400 1900 2415
rect 1950 2400 2050 2415
rect 2100 2400 2200 2415
rect 2250 2400 2350 2415
rect 0 -15 100 0
rect 150 -15 250 0
rect 300 -15 400 0
rect 450 -15 550 0
rect 600 -15 700 0
rect 750 -15 850 0
rect 900 -15 1000 0
rect 1050 -15 1150 0
rect 1200 -15 1300 0
rect 1350 -15 1450 0
rect 1500 -15 1600 0
rect 1650 -15 1750 0
rect 1800 -15 1900 0
rect 1950 -15 2050 0
rect 2100 -15 2200 0
rect 2250 -15 2350 0
<< locali >>
rect -95 2385 -5 2395
rect -95 15 -85 2385
rect -60 15 -40 2385
rect -15 15 -5 2385
rect -95 5 -5 15
rect 2355 2385 2445 2395
rect 2355 15 2365 2385
rect 2390 15 2410 2385
rect 2435 15 2445 2385
rect 2355 5 2445 15
<< end >>
