magic
tech sky130A
timestamp 1699558734
<< nwell >>
rect -120 2780 2470 4020
<< nmos >>
rect 0 1200 100 2400
rect 150 1200 250 2400
rect 300 1200 400 2400
rect 450 1200 550 2400
rect 600 1200 700 2400
rect 750 1200 850 2400
rect 900 1200 1000 2400
rect 1050 1200 1150 2400
rect 1200 1200 1300 2400
rect 1350 1200 1450 2400
rect 1500 1200 1600 2400
rect 1650 1200 1750 2400
rect 1800 1200 1900 2400
rect 1950 1200 2050 2400
rect 2100 1200 2200 2400
rect 2250 1200 2350 2400
<< pmos >>
rect 0 2800 100 4000
rect 150 2800 250 4000
rect 300 2800 400 4000
rect 530 2800 630 4000
rect 660 2800 760 4000
rect 790 2800 890 4000
rect 920 2800 1020 4000
rect 1050 2800 1150 4000
rect 1200 2800 1300 4000
rect 1330 2800 1430 4000
rect 1460 2800 1560 4000
rect 1590 2800 1690 4000
rect 1720 2800 1820 4000
rect 1950 2800 2050 4000
rect 2100 2800 2200 4000
rect 2250 2800 2350 4000
<< ndiff >>
rect -50 2385 0 2400
rect -50 1215 -40 2385
rect -15 1215 0 2385
rect -50 1200 0 1215
rect 100 2385 150 2400
rect 100 1215 115 2385
rect 135 1215 150 2385
rect 100 1200 150 1215
rect 250 2385 300 2400
rect 250 1215 265 2385
rect 285 1215 300 2385
rect 250 1200 300 1215
rect 400 2385 450 2400
rect 400 1215 415 2385
rect 435 1215 450 2385
rect 400 1200 450 1215
rect 550 2385 600 2400
rect 550 1215 565 2385
rect 585 1215 600 2385
rect 550 1200 600 1215
rect 700 2385 750 2400
rect 700 1215 715 2385
rect 735 1215 750 2385
rect 700 1200 750 1215
rect 850 2385 900 2400
rect 850 1215 865 2385
rect 885 1215 900 2385
rect 850 1200 900 1215
rect 1000 2385 1050 2400
rect 1000 1215 1015 2385
rect 1035 1215 1050 2385
rect 1000 1200 1050 1215
rect 1150 2385 1200 2400
rect 1150 1215 1165 2385
rect 1185 1215 1200 2385
rect 1150 1200 1200 1215
rect 1300 2385 1350 2400
rect 1300 1215 1315 2385
rect 1335 1215 1350 2385
rect 1300 1200 1350 1215
rect 1450 2385 1500 2400
rect 1450 1215 1465 2385
rect 1485 1215 1500 2385
rect 1450 1200 1500 1215
rect 1600 2385 1650 2400
rect 1600 1215 1615 2385
rect 1635 1215 1650 2385
rect 1600 1200 1650 1215
rect 1750 2385 1800 2400
rect 1750 1215 1765 2385
rect 1785 1215 1800 2385
rect 1750 1200 1800 1215
rect 1900 2385 1950 2400
rect 1900 1215 1915 2385
rect 1935 1215 1950 2385
rect 1900 1200 1950 1215
rect 2050 2385 2100 2400
rect 2050 1215 2065 2385
rect 2085 1215 2100 2385
rect 2050 1200 2100 1215
rect 2200 2385 2250 2400
rect 2200 1215 2215 2385
rect 2235 1215 2250 2385
rect 2200 1200 2250 1215
rect 2350 2385 2400 2400
rect 2350 1215 2365 2385
rect 2390 1215 2400 2385
rect 2350 1200 2400 1215
<< pdiff >>
rect -50 3985 0 4000
rect -50 2815 -40 3985
rect -15 2815 0 3985
rect -50 2800 0 2815
rect 100 3985 150 4000
rect 100 2815 115 3985
rect 135 2815 150 3985
rect 100 2800 150 2815
rect 250 3985 300 4000
rect 250 2815 265 3985
rect 285 2815 300 3985
rect 250 2800 300 2815
rect 400 3985 450 4000
rect 400 2815 415 3985
rect 435 2815 450 3985
rect 400 2800 450 2815
rect 480 3985 530 4000
rect 480 2815 495 3985
rect 515 2815 530 3985
rect 480 2800 530 2815
rect 630 2800 660 4000
rect 760 2800 790 4000
rect 890 2800 920 4000
rect 1020 2800 1050 4000
rect 1150 3985 1200 4000
rect 1150 2815 1165 3985
rect 1185 2815 1200 3985
rect 1150 2800 1200 2815
rect 1300 2800 1330 4000
rect 1430 2800 1460 4000
rect 1560 2800 1590 4000
rect 1690 2800 1720 4000
rect 1820 3985 1870 4000
rect 1820 2815 1835 3985
rect 1855 2815 1870 3985
rect 1820 2800 1870 2815
rect 1900 3985 1950 4000
rect 1900 2815 1915 3985
rect 1935 2815 1950 3985
rect 1900 2800 1950 2815
rect 2050 3985 2100 4000
rect 2050 2815 2065 3985
rect 2085 2815 2100 3985
rect 2050 2800 2100 2815
rect 2200 3985 2250 4000
rect 2200 2815 2215 3985
rect 2235 2815 2250 3985
rect 2200 2800 2250 2815
rect 2350 3985 2400 4000
rect 2350 2815 2365 3985
rect 2390 2815 2400 3985
rect 2350 2800 2400 2815
<< ndiffc >>
rect -40 1215 -15 2385
rect 115 1215 135 2385
rect 265 1215 285 2385
rect 415 1215 435 2385
rect 565 1215 585 2385
rect 715 1215 735 2385
rect 865 1215 885 2385
rect 1015 1215 1035 2385
rect 1165 1215 1185 2385
rect 1315 1215 1335 2385
rect 1465 1215 1485 2385
rect 1615 1215 1635 2385
rect 1765 1215 1785 2385
rect 1915 1215 1935 2385
rect 2065 1215 2085 2385
rect 2215 1215 2235 2385
rect 2365 1215 2390 2385
<< pdiffc >>
rect -40 2815 -15 3985
rect 115 2815 135 3985
rect 265 2815 285 3985
rect 415 2815 435 3985
rect 495 2815 515 3985
rect 1165 2815 1185 3985
rect 1835 2815 1855 3985
rect 1915 2815 1935 3985
rect 2065 2815 2085 3985
rect 2215 2815 2235 3985
rect 2365 2815 2390 3985
<< psubdiff >>
rect -100 2385 -50 2400
rect -100 1215 -85 2385
rect -60 1215 -50 2385
rect -100 1200 -50 1215
rect 2400 2385 2450 2400
rect 2400 1215 2410 2385
rect 2435 1215 2450 2385
rect 2400 1200 2450 1215
<< nsubdiff >>
rect -100 3985 -50 4000
rect -100 2815 -85 3985
rect -60 2815 -50 3985
rect -100 2800 -50 2815
rect 2400 3985 2450 4000
rect 2400 2815 2410 3985
rect 2435 2815 2450 3985
rect 2400 2800 2450 2815
<< psubdiffcont >>
rect -85 1215 -60 2385
rect 2410 1215 2435 2385
<< nsubdiffcont >>
rect -85 2815 -60 3985
rect 2410 2815 2435 3985
<< poly >>
rect 0 4000 100 4015
rect 150 4000 250 4015
rect 300 4000 400 4015
rect 530 4000 630 4015
rect 660 4000 760 4015
rect 790 4000 890 4015
rect 920 4000 1020 4015
rect 1050 4000 1150 4015
rect 1200 4000 1300 4015
rect 1330 4000 1430 4015
rect 1460 4000 1560 4015
rect 1590 4000 1690 4015
rect 1720 4000 1820 4015
rect 1950 4000 2050 4015
rect 2100 4000 2200 4015
rect 2250 4000 2350 4015
rect 0 2785 100 2800
rect 150 2785 250 2800
rect 300 2785 400 2800
rect 530 2785 630 2800
rect 660 2785 760 2800
rect 790 2785 890 2800
rect 920 2785 1020 2800
rect 1050 2785 1150 2800
rect 1200 2785 1300 2800
rect 1330 2785 1430 2800
rect 1460 2785 1560 2800
rect 1590 2785 1690 2800
rect 1720 2785 1820 2800
rect 1950 2785 2050 2800
rect 2100 2785 2200 2800
rect 2250 2785 2350 2800
rect 0 2400 100 2415
rect 150 2400 250 2415
rect 300 2400 400 2415
rect 450 2400 550 2415
rect 600 2400 700 2415
rect 750 2400 850 2415
rect 900 2400 1000 2415
rect 1050 2400 1150 2415
rect 1200 2400 1300 2415
rect 1350 2400 1450 2415
rect 1500 2400 1600 2415
rect 1650 2400 1750 2415
rect 1800 2400 1900 2415
rect 1950 2400 2050 2415
rect 2100 2400 2200 2415
rect 2250 2400 2350 2415
rect 0 1185 100 1200
rect 150 1185 250 1200
rect 300 1160 400 1200
rect 450 1160 550 1200
rect 600 1160 700 1200
rect 750 1160 850 1200
rect 900 1160 1000 1200
rect 1050 1185 1150 1200
rect 1200 1185 1300 1200
rect 1350 1160 1450 1200
rect 1500 1160 1600 1200
rect 1650 1160 1750 1200
rect 1800 1160 1900 1200
rect 1950 1160 2050 1200
rect 2100 1185 2200 1200
rect 2250 1185 2350 1200
rect 300 1145 2050 1160
<< locali >>
rect -95 3985 -5 3995
rect -95 2815 -85 3985
rect -60 2815 -40 3985
rect -15 2815 -5 3985
rect -95 2805 -5 2815
rect 105 3985 145 3995
rect 105 2815 115 3985
rect 135 2815 145 3985
rect 105 2805 145 2815
rect 255 3985 295 3995
rect 255 2815 265 3985
rect 285 2815 295 3985
rect 255 2805 295 2815
rect 405 3985 445 3995
rect 405 2815 415 3985
rect 435 2815 445 3985
rect 405 2805 445 2815
rect 485 3985 525 3995
rect 485 2815 495 3985
rect 515 2815 525 3985
rect 485 2805 525 2815
rect 1155 3985 1195 3995
rect 1155 2815 1165 3985
rect 1185 2815 1195 3985
rect 1155 2805 1195 2815
rect 1825 3985 1865 3995
rect 1825 2815 1835 3985
rect 1855 2815 1865 3985
rect 1825 2805 1865 2815
rect 1905 3985 1945 3995
rect 1905 2815 1915 3985
rect 1935 2815 1945 3985
rect 1905 2805 1945 2815
rect 2055 3985 2095 3995
rect 2055 2815 2065 3985
rect 2085 2815 2095 3985
rect 2055 2805 2095 2815
rect 2205 3985 2245 3995
rect 2205 2815 2215 3985
rect 2235 2815 2245 3985
rect 2205 2805 2245 2815
rect 2355 3985 2445 3995
rect 2355 2815 2365 3985
rect 2390 2815 2410 3985
rect 2435 2815 2445 3985
rect 2355 2805 2445 2815
rect 555 2415 1795 2435
rect -95 2385 -5 2395
rect -95 1215 -85 2385
rect -60 1215 -40 2385
rect -15 1215 -5 2385
rect -95 1205 -5 1215
rect 105 2385 145 2395
rect 105 1215 115 2385
rect 135 1215 145 2385
rect 105 1205 145 1215
rect 255 2385 295 2395
rect 255 1215 265 2385
rect 285 1215 295 2385
rect 255 1205 295 1215
rect 405 2385 445 2395
rect 405 1215 415 2385
rect 435 1215 445 2385
rect 405 1185 445 1215
rect 555 2385 595 2415
rect 555 1215 565 2385
rect 585 1215 595 2385
rect 555 1205 595 1215
rect 705 2385 745 2395
rect 705 1215 715 2385
rect 735 1215 745 2385
rect 705 1185 745 1215
rect 855 2385 895 2415
rect 855 1215 865 2385
rect 885 1215 895 2385
rect 855 1205 895 1215
rect 1005 2385 1045 2395
rect 1005 1215 1015 2385
rect 1035 1215 1045 2385
rect 1005 1185 1045 1215
rect 1155 2385 1195 2395
rect 1155 1215 1165 2385
rect 1185 1215 1195 2385
rect 1155 1205 1195 1215
rect 1305 2385 1345 2395
rect 1305 1215 1315 2385
rect 1335 1215 1345 2385
rect 1305 1185 1345 1215
rect 1455 2385 1495 2415
rect 1455 1215 1465 2385
rect 1485 1215 1495 2385
rect 1455 1205 1495 1215
rect 1605 2385 1645 2395
rect 1605 1215 1615 2385
rect 1635 1215 1645 2385
rect 1605 1185 1645 1215
rect 1755 2385 1795 2415
rect 1755 1215 1765 2385
rect 1785 1215 1795 2385
rect 1755 1205 1795 1215
rect 1905 2385 1945 2395
rect 1905 1215 1915 2385
rect 1935 1215 1945 2385
rect 1905 1185 1945 1215
rect 2055 2385 2095 2395
rect 2055 1215 2065 2385
rect 2085 1215 2095 2385
rect 2055 1205 2095 1215
rect 2205 2385 2245 2395
rect 2205 1215 2215 2385
rect 2235 1215 2245 2385
rect 2205 1205 2245 1215
rect 2355 2385 2445 2395
rect 2355 1215 2365 2385
rect 2390 1215 2410 2385
rect 2435 1215 2445 2385
rect 2355 1205 2445 1215
rect 405 1165 1945 1185
<< end >>
