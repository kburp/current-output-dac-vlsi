magic
tech sky130A
timestamp 1699588500
<< nwell >>
rect 2314 164 2602 2640
<< nmos >>
rect 0 200 100 2600
rect 150 200 250 2600
rect 300 200 400 2600
rect 450 200 550 2600
rect 600 200 700 2600
rect 750 200 850 2600
rect 900 200 1000 2600
rect 1050 200 1150 2600
rect 1200 200 1300 2600
rect 1350 200 1450 2600
rect 1500 200 1600 2600
rect 1650 200 1750 2600
rect 1800 200 1900 2600
rect 1950 200 2050 2600
rect 2100 200 2200 2600
rect 0 -2400 100 0
rect 150 -2400 250 0
rect 300 -2400 400 0
rect 450 -2400 550 0
rect 600 -2400 700 0
rect 750 -2400 850 0
rect 900 -2400 1000 0
rect 1050 -2400 1150 0
rect 1200 -2400 1300 0
rect 1350 -2400 1450 0
rect 1500 -2400 1600 0
rect 1650 -2400 1750 0
rect 1800 -2400 1900 0
rect 1950 -2400 2050 0
rect 2100 -2400 2200 0
rect 2250 -2400 2350 0
rect 2400 -2400 2500 0
<< pmos >>
rect 2384 200 2484 2600
<< ndiff >>
rect -50 2578 0 2600
rect -50 222 -34 2578
rect -16 222 0 2578
rect -50 200 0 222
rect 100 2578 150 2600
rect 100 222 116 2578
rect 134 222 150 2578
rect 100 200 150 222
rect 250 2578 300 2600
rect 250 222 266 2578
rect 284 222 300 2578
rect 250 200 300 222
rect 400 2578 450 2600
rect 400 222 416 2578
rect 434 222 450 2578
rect 400 200 450 222
rect 550 2578 600 2600
rect 550 222 566 2578
rect 584 222 600 2578
rect 550 200 600 222
rect 700 2578 750 2600
rect 700 222 716 2578
rect 734 222 750 2578
rect 700 200 750 222
rect 850 2578 900 2600
rect 850 222 866 2578
rect 884 222 900 2578
rect 850 200 900 222
rect 1000 2578 1050 2600
rect 1000 222 1016 2578
rect 1034 222 1050 2578
rect 1000 200 1050 222
rect 1150 2578 1200 2600
rect 1150 222 1166 2578
rect 1184 222 1200 2578
rect 1150 200 1200 222
rect 1300 2578 1350 2600
rect 1300 222 1316 2578
rect 1334 222 1350 2578
rect 1300 200 1350 222
rect 1450 2578 1500 2600
rect 1450 222 1466 2578
rect 1484 222 1500 2578
rect 1450 200 1500 222
rect 1600 2578 1650 2600
rect 1600 222 1616 2578
rect 1634 222 1650 2578
rect 1600 200 1650 222
rect 1750 2578 1800 2600
rect 1750 222 1766 2578
rect 1784 222 1800 2578
rect 1750 200 1800 222
rect 1900 2578 1950 2600
rect 1900 222 1916 2578
rect 1934 222 1950 2578
rect 1900 200 1950 222
rect 2050 2578 2100 2600
rect 2050 222 2066 2578
rect 2084 222 2100 2578
rect 2050 200 2100 222
rect 2200 2578 2250 2600
rect 2200 222 2216 2578
rect 2234 222 2250 2578
rect 2200 200 2250 222
rect -50 -22 0 0
rect -50 -2378 -34 -22
rect -16 -2378 0 -22
rect -50 -2400 0 -2378
rect 100 -22 150 0
rect 100 -2378 116 -22
rect 134 -2378 150 -22
rect 100 -2400 150 -2378
rect 250 -22 300 0
rect 250 -2378 266 -22
rect 284 -2378 300 -22
rect 250 -2400 300 -2378
rect 400 -22 450 0
rect 400 -2378 416 -22
rect 434 -2378 450 -22
rect 400 -2400 450 -2378
rect 550 -22 600 0
rect 550 -2378 566 -22
rect 584 -2378 600 -22
rect 550 -2400 600 -2378
rect 700 -22 750 0
rect 700 -2378 716 -22
rect 734 -2378 750 -22
rect 700 -2400 750 -2378
rect 850 -22 900 0
rect 850 -2378 866 -22
rect 884 -2378 900 -22
rect 850 -2400 900 -2378
rect 1000 -22 1050 0
rect 1000 -2378 1016 -22
rect 1034 -2378 1050 -22
rect 1000 -2400 1050 -2378
rect 1150 -22 1200 0
rect 1150 -2378 1166 -22
rect 1184 -2378 1200 -22
rect 1150 -2400 1200 -2378
rect 1300 -22 1350 0
rect 1300 -2378 1316 -22
rect 1334 -2378 1350 -22
rect 1300 -2400 1350 -2378
rect 1450 -22 1500 0
rect 1450 -2378 1466 -22
rect 1484 -2378 1500 -22
rect 1450 -2400 1500 -2378
rect 1600 -22 1650 0
rect 1600 -2378 1616 -22
rect 1634 -2378 1650 -22
rect 1600 -2400 1650 -2378
rect 1750 -22 1800 0
rect 1750 -2378 1766 -22
rect 1784 -2378 1800 -22
rect 1750 -2400 1800 -2378
rect 1900 -22 1950 0
rect 1900 -2378 1916 -22
rect 1934 -2378 1950 -22
rect 1900 -2400 1950 -2378
rect 2050 -22 2100 0
rect 2050 -2378 2066 -22
rect 2084 -2378 2100 -22
rect 2050 -2400 2100 -2378
rect 2200 -22 2250 0
rect 2200 -2378 2216 -22
rect 2234 -2378 2250 -22
rect 2200 -2400 2250 -2378
rect 2350 -22 2400 0
rect 2350 -2378 2366 -22
rect 2384 -2378 2400 -22
rect 2350 -2400 2400 -2378
rect 2500 -22 2550 0
rect 2500 -2378 2516 -22
rect 2534 -2378 2550 -22
rect 2500 -2400 2550 -2378
<< pdiff >>
rect 2334 2578 2384 2600
rect 2334 222 2350 2578
rect 2368 222 2384 2578
rect 2334 200 2384 222
rect 2484 2578 2534 2600
rect 2484 222 2500 2578
rect 2518 222 2534 2578
rect 2484 200 2534 222
<< ndiffc >>
rect -34 222 -16 2578
rect 116 222 134 2578
rect 266 222 284 2578
rect 416 222 434 2578
rect 566 222 584 2578
rect 716 222 734 2578
rect 866 222 884 2578
rect 1016 222 1034 2578
rect 1166 222 1184 2578
rect 1316 222 1334 2578
rect 1466 222 1484 2578
rect 1616 222 1634 2578
rect 1766 222 1784 2578
rect 1916 222 1934 2578
rect 2066 222 2084 2578
rect 2216 222 2234 2578
rect -34 -2378 -16 -22
rect 116 -2378 134 -22
rect 266 -2378 284 -22
rect 416 -2378 434 -22
rect 566 -2378 584 -22
rect 716 -2378 734 -22
rect 866 -2378 884 -22
rect 1016 -2378 1034 -22
rect 1166 -2378 1184 -22
rect 1316 -2378 1334 -22
rect 1466 -2378 1484 -22
rect 1616 -2378 1634 -22
rect 1766 -2378 1784 -22
rect 1916 -2378 1934 -22
rect 2066 -2378 2084 -22
rect 2216 -2378 2234 -22
rect 2366 -2378 2384 -22
rect 2516 -2378 2534 -22
<< pdiffc >>
rect 2350 222 2368 2578
rect 2500 222 2518 2578
<< psubdiff >>
rect -100 2577 -50 2600
rect -100 237 -84 2577
rect -66 237 -50 2577
rect -100 200 -50 237
rect 2250 2576 2300 2600
rect 2250 220 2267 2576
rect 2287 220 2300 2576
rect 2250 200 2300 220
rect -100 -21 -50 0
rect -100 -2377 -81 -21
rect -63 -2377 -50 -21
rect -100 -2400 -50 -2377
rect 2550 -29 2600 0
rect 2550 -2379 2568 -29
rect 2585 -2379 2600 -29
rect 2550 -2400 2600 -2379
<< nsubdiff >>
rect 2534 2577 2584 2600
rect 2534 221 2550 2577
rect 2570 221 2584 2577
rect 2534 200 2584 221
<< psubdiffcont >>
rect -84 237 -66 2577
rect 2267 220 2287 2576
rect -81 -2377 -63 -21
rect 2568 -2379 2585 -29
<< nsubdiffcont >>
rect 2550 221 2570 2577
<< poly >>
rect 0 2600 100 2615
rect 150 2600 250 2615
rect 300 2600 400 2615
rect 450 2600 550 2615
rect 600 2600 700 2615
rect 750 2600 850 2615
rect 900 2600 1000 2615
rect 1050 2600 1150 2615
rect 1200 2600 1300 2615
rect 1350 2600 1450 2615
rect 1500 2600 1600 2615
rect 1650 2600 1750 2615
rect 1800 2600 1900 2615
rect 1950 2600 2050 2615
rect 2100 2600 2200 2615
rect 2384 2600 2484 2615
rect 0 160 100 200
rect 0 134 25 160
rect 55 134 100 160
rect 0 0 100 134
rect 150 185 250 200
rect 300 185 400 200
rect 450 185 550 200
rect 600 185 700 200
rect 750 185 850 200
rect 900 185 1000 200
rect 1050 185 1150 200
rect 1200 185 1300 200
rect 1350 185 1450 200
rect 1500 185 1600 200
rect 1650 185 1750 200
rect 1800 185 1900 200
rect 1950 185 2050 200
rect 150 170 700 185
rect 1050 170 1900 185
rect 2100 180 2200 200
rect 150 30 250 170
rect 1050 65 1150 170
rect 2100 160 2110 180
rect 2190 160 2200 180
rect 2100 155 2200 160
rect 2384 174 2484 200
rect 2384 155 2407 174
rect 2453 155 2484 174
rect 2384 143 2484 155
rect 1451 125 1498 128
rect 2384 125 2400 143
rect 1451 121 2400 125
rect 1451 102 1460 121
rect 1490 110 2400 121
rect 1490 102 1498 110
rect 1451 94 1498 102
rect 600 50 1150 65
rect 2335 70 2545 85
rect 2335 55 2350 70
rect 600 30 700 50
rect 150 15 700 30
rect 1050 30 1150 50
rect 1800 40 2350 55
rect 1800 30 1900 40
rect 1050 15 1900 30
rect 150 0 250 15
rect 300 0 400 15
rect 450 0 550 15
rect 600 0 700 15
rect 750 0 850 15
rect 900 0 1000 15
rect 1050 0 1150 15
rect 1200 0 1300 15
rect 1350 0 1450 15
rect 1500 0 1600 15
rect 1650 0 1750 15
rect 1800 0 1900 15
rect 1950 0 2050 15
rect 2100 0 2200 15
rect 2250 0 2350 40
rect 2400 37 2500 45
rect 2400 20 2430 37
rect 2465 20 2500 37
rect 2400 0 2500 20
rect 0 -2415 100 -2400
rect 150 -2415 250 -2400
rect 300 -2415 400 -2400
rect 450 -2415 550 -2400
rect 600 -2415 700 -2400
rect 750 -2415 850 -2400
rect 900 -2415 1000 -2400
rect 1050 -2415 1150 -2400
rect 1200 -2415 1300 -2400
rect 1350 -2415 1450 -2400
rect 1500 -2415 1600 -2400
rect 1650 -2415 1750 -2400
rect 1800 -2415 1900 -2400
rect 1950 -2415 2050 -2400
rect 2100 -2415 2200 -2400
rect 2250 -2415 2350 -2400
rect 2400 -2415 2500 -2400
<< polycont >>
rect 25 134 55 160
rect 2110 160 2190 180
rect 2407 155 2453 174
rect 1460 102 1490 121
rect 2430 20 2465 37
<< locali >>
rect 260 2642 1040 2659
rect -90 2577 -60 2589
rect -90 237 -84 2577
rect -66 237 -60 2577
rect -90 209 -60 237
rect -40 2578 -10 2590
rect -40 222 -34 2578
rect -16 222 -10 2578
rect -40 170 -10 222
rect 110 2578 140 2590
rect 110 222 116 2578
rect 134 222 140 2578
rect 110 192 140 222
rect 260 2578 290 2642
rect 260 222 266 2578
rect 284 222 290 2578
rect 260 210 290 222
rect 410 2607 740 2624
rect 410 2578 440 2607
rect 410 222 416 2578
rect 434 222 440 2578
rect 410 192 440 222
rect 110 175 440 192
rect 560 2578 590 2590
rect 560 222 566 2578
rect 584 222 590 2578
rect -40 160 70 170
rect -40 150 25 160
rect 10 134 25 150
rect 55 134 70 160
rect 10 120 70 134
rect 560 122 590 222
rect 710 2578 740 2607
rect 710 222 716 2578
rect 734 222 740 2578
rect 710 199 740 222
rect 860 2578 890 2590
rect 860 222 866 2578
rect 884 222 890 2578
rect 860 210 890 222
rect 1010 2578 1040 2642
rect 1010 222 1016 2578
rect 1034 222 1040 2578
rect 1010 193 1040 222
rect 1160 2613 1940 2630
rect 1160 2608 1640 2613
rect 1160 2578 1190 2608
rect 1160 222 1166 2578
rect 1184 222 1190 2578
rect 1160 210 1190 222
rect 1310 2578 1340 2590
rect 1310 222 1316 2578
rect 1334 222 1340 2578
rect 1310 193 1340 222
rect 1010 176 1340 193
rect 1460 2578 1490 2590
rect 1460 222 1466 2578
rect 1484 222 1490 2578
rect 1460 128 1490 222
rect 1610 2578 1640 2608
rect 1610 222 1616 2578
rect 1634 222 1640 2578
rect 1610 210 1640 222
rect 1760 2578 1790 2590
rect 1760 222 1766 2578
rect 1784 222 1790 2578
rect 1451 122 1498 128
rect 560 121 1498 122
rect 560 102 1460 121
rect 1490 102 1498 121
rect 560 101 1498 102
rect 1451 94 1498 101
rect -102 13 290 30
rect -87 -21 -57 -7
rect -87 -2377 -81 -21
rect -63 -2377 -57 -21
rect -87 -2387 -57 -2377
rect -40 -22 -10 -10
rect -40 -2378 -34 -22
rect -16 -2378 -10 -22
rect -40 -2390 -10 -2378
rect 110 -22 140 -10
rect 110 -2378 116 -22
rect 134 -2378 140 -22
rect 110 -2418 140 -2378
rect 260 -22 290 13
rect 560 8 1340 25
rect 260 -2378 266 -22
rect 284 -2378 290 -22
rect 260 -2390 290 -2378
rect 410 -22 440 -10
rect 410 -2378 416 -22
rect 434 -2378 440 -22
rect 410 -2418 440 -2378
rect 560 -22 590 8
rect 560 -2378 566 -22
rect 584 -2378 590 -22
rect 560 -2390 590 -2378
rect 710 -22 740 -10
rect 710 -2378 716 -22
rect 734 -2378 740 -22
rect 710 -2418 740 -2378
rect 860 -22 890 -10
rect 860 -2378 866 -22
rect 884 -2378 890 -22
rect 860 -2390 890 -2378
rect 1010 -22 1040 8
rect 1010 -2378 1016 -22
rect 1034 -2378 1040 -22
rect 1010 -2390 1040 -2378
rect 1160 -22 1190 -10
rect 1160 -2378 1166 -22
rect 1184 -2378 1190 -22
rect 110 -2435 740 -2418
rect 1160 -2408 1190 -2378
rect 1310 -22 1340 8
rect 1310 -2378 1316 -22
rect 1334 -2378 1340 -22
rect 1310 -2390 1340 -2378
rect 1460 -22 1490 94
rect 1760 33 1790 222
rect 1910 2578 1940 2613
rect 1910 222 1916 2578
rect 1934 222 1940 2578
rect 1910 210 1940 222
rect 2060 2578 2090 2590
rect 2060 222 2066 2578
rect 2084 222 2090 2578
rect 2060 185 2090 222
rect 2210 2578 2240 2590
rect 2210 222 2216 2578
rect 2234 222 2240 2578
rect 2210 210 2240 222
rect 2261 2576 2291 2591
rect 2261 220 2267 2576
rect 2287 220 2291 2576
rect 2261 211 2291 220
rect 2344 2578 2374 2590
rect 2344 222 2350 2578
rect 2368 222 2374 2578
rect 2060 180 2200 185
rect 2060 160 2110 180
rect 2190 160 2200 180
rect 2060 155 2200 160
rect 2344 154 2374 222
rect 2494 2578 2524 2590
rect 2494 222 2500 2578
rect 2518 222 2524 2578
rect 2494 210 2524 222
rect 2545 2577 2575 2596
rect 2545 221 2550 2577
rect 2570 221 2575 2577
rect 2545 208 2575 221
rect 2394 174 2466 179
rect 2394 163 2407 174
rect 2391 155 2407 163
rect 2453 155 2466 174
rect 2391 154 2466 155
rect 2344 146 2466 154
rect 2344 128 2408 146
rect 2360 127 2408 128
rect 1760 16 2240 33
rect 1460 -2378 1466 -22
rect 1484 -2378 1490 -22
rect 1460 -2390 1490 -2378
rect 1610 -22 1640 -10
rect 1610 -2378 1616 -22
rect 1634 -2378 1640 -22
rect 1610 -2408 1640 -2378
rect 1760 -22 1790 16
rect 1760 -2378 1766 -22
rect 1784 -2378 1790 -22
rect 1760 -2390 1790 -2378
rect 1910 -22 1940 -10
rect 1910 -2378 1916 -22
rect 1934 -2378 1940 -22
rect 1910 -2408 1940 -2378
rect 2060 -22 2090 -10
rect 2060 -2378 2066 -22
rect 2084 -2378 2090 -22
rect 2060 -2390 2090 -2378
rect 2210 -22 2240 16
rect 2210 -2378 2216 -22
rect 2234 -2378 2240 -22
rect 2210 -2390 2240 -2378
rect 2360 -22 2390 127
rect 2422 37 2477 45
rect 2422 20 2430 37
rect 2465 20 2541 37
rect 2422 15 2541 20
rect 2422 5 2475 15
rect 2509 -18 2541 15
rect 2360 -2378 2366 -22
rect 2384 -2378 2390 -22
rect 2360 -2390 2390 -2378
rect 2510 -22 2540 -18
rect 2510 -2378 2516 -22
rect 2534 -2378 2540 -22
rect 2510 -2390 2540 -2378
rect 2561 -29 2590 -17
rect 2561 -2379 2568 -29
rect 2585 -2379 2590 -29
rect 2561 -2388 2590 -2379
rect 1160 -2426 1940 -2408
<< viali >>
rect -84 237 -66 2577
rect -34 222 -16 2578
rect 866 222 884 2578
rect -34 -2378 -16 -22
rect 866 -2378 884 -22
rect 2066 222 2084 2578
rect 2216 222 2234 2578
rect 2267 220 2287 2576
rect 2500 222 2518 2578
rect 2550 221 2570 2577
rect 2066 -2378 2084 -22
rect 2516 -2378 2534 -22
rect 2568 -2379 2585 -29
<< metal1 >>
rect -100 2577 -54 2600
rect -100 237 -87 2577
rect -61 237 -54 2577
rect -100 200 -54 237
rect -40 2578 -10 2585
rect -40 222 -38 2578
rect -12 222 -10 2578
rect -40 210 -10 222
rect 860 2578 890 2585
rect 860 222 862 2578
rect 888 222 890 2578
rect 860 210 890 222
rect 2060 2578 2090 2585
rect 2060 222 2062 2578
rect 2088 222 2090 2578
rect 2060 210 2090 222
rect 2210 2578 2240 2585
rect 2210 222 2212 2578
rect 2238 222 2240 2578
rect 2210 210 2240 222
rect 2254 2577 2300 2600
rect 2254 220 2258 2577
rect 2294 220 2300 2577
rect 2254 200 2300 220
rect 2484 2578 2584 2600
rect 2484 222 2496 2578
rect 2522 2577 2584 2578
rect 2522 222 2547 2577
rect 2484 221 2547 222
rect 2573 221 2584 2577
rect 2484 200 2584 221
rect -41 -22 -9 -9
rect -41 -2378 -38 -22
rect -12 -2378 -9 -22
rect -41 -2391 -9 -2378
rect 859 -22 891 -9
rect 859 -2378 862 -22
rect 888 -2378 891 -22
rect 859 -2391 891 -2378
rect 2059 -22 2091 -9
rect 2059 -2378 2062 -22
rect 2088 -2378 2091 -22
rect 2059 -2391 2091 -2378
rect 2509 -22 2541 -9
rect 2509 -2378 2512 -22
rect 2538 -2378 2541 -22
rect 2509 -2391 2541 -2378
rect 2555 -29 2600 0
rect 2555 -2379 2562 -29
rect 2588 -2379 2600 -29
rect 2555 -2400 2600 -2379
<< via1 >>
rect -87 237 -84 2577
rect -84 237 -66 2577
rect -66 237 -61 2577
rect -38 222 -34 2578
rect -34 222 -16 2578
rect -16 222 -12 2578
rect 862 222 866 2578
rect 866 222 884 2578
rect 884 222 888 2578
rect 2062 222 2066 2578
rect 2066 222 2084 2578
rect 2084 222 2088 2578
rect 2212 222 2216 2578
rect 2216 222 2234 2578
rect 2234 222 2238 2578
rect 2258 2576 2294 2577
rect 2258 220 2267 2576
rect 2267 220 2287 2576
rect 2287 220 2294 2576
rect 2496 222 2500 2578
rect 2500 222 2518 2578
rect 2518 222 2522 2578
rect 2547 221 2550 2577
rect 2550 221 2570 2577
rect 2570 221 2573 2577
rect -38 -2378 -34 -22
rect -34 -2378 -16 -22
rect -16 -2378 -12 -22
rect 862 -2378 866 -22
rect 866 -2378 884 -22
rect 884 -2378 888 -22
rect 2062 -2378 2066 -22
rect 2066 -2378 2084 -22
rect 2084 -2378 2088 -22
rect 2512 -2378 2516 -22
rect 2516 -2378 2534 -22
rect 2534 -2378 2538 -22
rect 2562 -2379 2568 -29
rect 2568 -2379 2585 -29
rect 2585 -2379 2588 -29
<< metal2 >>
rect -100 2578 2300 2600
rect -100 2577 -38 2578
rect -100 237 -87 2577
rect -61 237 -38 2577
rect -100 222 -38 237
rect -12 222 862 2578
rect 888 222 2062 2578
rect 2088 222 2212 2578
rect 2238 2577 2300 2578
rect 2238 222 2258 2577
rect -100 220 2258 222
rect 2294 220 2300 2577
rect -100 202 2300 220
rect -101 0 2300 202
rect 2328 2578 2586 2599
rect 2328 222 2496 2578
rect 2522 2577 2586 2578
rect 2522 222 2547 2577
rect 2328 221 2547 222
rect 2573 221 2586 2577
rect 2328 198 2586 221
rect -101 -22 2602 0
rect -101 -2378 -38 -22
rect -12 -2378 862 -22
rect 888 -2378 2062 -22
rect 2088 -2378 2512 -22
rect 2538 -29 2602 -22
rect 2538 -2378 2562 -29
rect -101 -2379 2562 -2378
rect 2588 -2379 2602 -29
rect -101 -2400 2602 -2379
<< labels >>
rlabel poly 2545 77 2545 77 3 Vgate
rlabel locali -102 22 -102 22 7 Idac
rlabel metal2 -101 36 -101 36 7 VN
rlabel metal2 2586 201 2586 201 3 VP
rlabel poly 2149 -2415 2149 -2415 5 b3
rlabel poly 2000 -2415 2000 -2415 5 b4
rlabel poly 1999 2615 1999 2615 1 b2
rlabel poly 952 2615 952 2615 1 b1
rlabel poly 801 2615 801 2615 1 b0
rlabel poly 955 -2415 955 -2415 5 b5
rlabel poly 794 -2415 794 -2415 5 b6
<< end >>
