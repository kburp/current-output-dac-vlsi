magic
tech sky130A
timestamp 1699636225
<< nwell >>
rect -120 2490 2470 3730
<< nmos >>
rect 0 1200 100 2400
rect 150 1200 250 2400
rect 300 1200 400 2400
rect 450 1200 550 2400
rect 600 1200 700 2400
rect 750 1200 850 2400
rect 900 1200 1000 2400
rect 1050 1200 1150 2400
rect 1200 1200 1300 2400
rect 1350 1200 1450 2400
rect 1500 1200 1600 2400
rect 1650 1200 1750 2400
rect 1800 1200 1900 2400
rect 1950 1200 2050 2400
rect 2100 1200 2200 2400
rect 2250 1200 2350 2400
<< pmos >>
rect 0 2510 100 3710
rect 150 2510 250 3710
rect 300 2510 400 3710
rect 530 2510 630 3710
rect 660 2510 760 3710
rect 790 2510 890 3710
rect 920 2510 1020 3710
rect 1050 2510 1150 3710
rect 1200 2510 1300 3710
rect 1330 2510 1430 3710
rect 1460 2510 1560 3710
rect 1590 2510 1690 3710
rect 1720 2510 1820 3710
rect 1950 2510 2050 3710
rect 2100 2510 2200 3710
rect 2250 2510 2350 3710
<< ndiff >>
rect -50 2385 0 2400
rect -50 1215 -40 2385
rect -15 1215 0 2385
rect -50 1200 0 1215
rect 100 2385 150 2400
rect 100 1215 115 2385
rect 135 1215 150 2385
rect 100 1200 150 1215
rect 250 2385 300 2400
rect 250 1215 265 2385
rect 285 1215 300 2385
rect 250 1200 300 1215
rect 400 2385 450 2400
rect 400 1215 415 2385
rect 435 1215 450 2385
rect 400 1200 450 1215
rect 550 2385 600 2400
rect 550 1215 565 2385
rect 585 1215 600 2385
rect 550 1200 600 1215
rect 700 2385 750 2400
rect 700 1215 715 2385
rect 735 1215 750 2385
rect 700 1200 750 1215
rect 850 2385 900 2400
rect 850 1215 865 2385
rect 885 1215 900 2385
rect 850 1200 900 1215
rect 1000 2385 1050 2400
rect 1000 1215 1015 2385
rect 1035 1215 1050 2385
rect 1000 1200 1050 1215
rect 1150 2385 1200 2400
rect 1150 1215 1165 2385
rect 1185 1215 1200 2385
rect 1150 1200 1200 1215
rect 1300 2385 1350 2400
rect 1300 1215 1315 2385
rect 1335 1215 1350 2385
rect 1300 1200 1350 1215
rect 1450 2385 1500 2400
rect 1450 1215 1465 2385
rect 1485 1215 1500 2385
rect 1450 1200 1500 1215
rect 1600 2385 1650 2400
rect 1600 1215 1615 2385
rect 1635 1215 1650 2385
rect 1600 1200 1650 1215
rect 1750 2385 1800 2400
rect 1750 1215 1765 2385
rect 1785 1215 1800 2385
rect 1750 1200 1800 1215
rect 1900 2385 1950 2400
rect 1900 1215 1915 2385
rect 1935 1215 1950 2385
rect 1900 1200 1950 1215
rect 2050 2385 2100 2400
rect 2050 1215 2065 2385
rect 2085 1215 2100 2385
rect 2050 1200 2100 1215
rect 2200 2385 2250 2400
rect 2200 1215 2215 2385
rect 2235 1215 2250 2385
rect 2200 1200 2250 1215
rect 2350 2385 2400 2400
rect 2350 1215 2365 2385
rect 2390 1215 2400 2385
rect 2350 1200 2400 1215
<< pdiff >>
rect -50 3695 0 3710
rect -50 2525 -40 3695
rect -15 2525 0 3695
rect -50 2510 0 2525
rect 100 3695 150 3710
rect 100 2525 115 3695
rect 135 2525 150 3695
rect 100 2510 150 2525
rect 250 3695 300 3710
rect 250 2525 265 3695
rect 285 2525 300 3695
rect 250 2510 300 2525
rect 400 3695 450 3710
rect 400 2525 415 3695
rect 435 2525 450 3695
rect 400 2510 450 2525
rect 480 3695 530 3710
rect 480 2525 495 3695
rect 515 2525 530 3695
rect 480 2510 530 2525
rect 630 2510 660 3710
rect 760 2510 790 3710
rect 890 2510 920 3710
rect 1020 2510 1050 3710
rect 1150 3695 1200 3710
rect 1150 2525 1165 3695
rect 1185 2525 1200 3695
rect 1150 2510 1200 2525
rect 1300 2510 1330 3710
rect 1430 2510 1460 3710
rect 1560 2510 1590 3710
rect 1690 2510 1720 3710
rect 1820 3695 1870 3710
rect 1820 2525 1835 3695
rect 1855 2525 1870 3695
rect 1820 2510 1870 2525
rect 1900 3695 1950 3710
rect 1900 2525 1915 3695
rect 1935 2525 1950 3695
rect 1900 2510 1950 2525
rect 2050 3695 2100 3710
rect 2050 2525 2065 3695
rect 2085 2525 2100 3695
rect 2050 2510 2100 2525
rect 2200 3695 2250 3710
rect 2200 2525 2215 3695
rect 2235 2525 2250 3695
rect 2200 2510 2250 2525
rect 2350 3695 2400 3710
rect 2350 2525 2365 3695
rect 2390 2525 2400 3695
rect 2350 2510 2400 2525
<< ndiffc >>
rect -40 1215 -15 2385
rect 115 1215 135 2385
rect 265 1215 285 2385
rect 415 1215 435 2385
rect 565 1215 585 2385
rect 715 1215 735 2385
rect 865 1215 885 2385
rect 1015 1215 1035 2385
rect 1165 1215 1185 2385
rect 1315 1215 1335 2385
rect 1465 1215 1485 2385
rect 1615 1215 1635 2385
rect 1765 1215 1785 2385
rect 1915 1215 1935 2385
rect 2065 1215 2085 2385
rect 2215 1215 2235 2385
rect 2365 1215 2390 2385
<< pdiffc >>
rect -40 2525 -15 3695
rect 115 2525 135 3695
rect 265 2525 285 3695
rect 415 2525 435 3695
rect 495 2525 515 3695
rect 1165 2525 1185 3695
rect 1835 2525 1855 3695
rect 1915 2525 1935 3695
rect 2065 2525 2085 3695
rect 2215 2525 2235 3695
rect 2365 2525 2390 3695
<< psubdiff >>
rect -100 2385 -50 2400
rect -100 1215 -85 2385
rect -60 1215 -50 2385
rect -100 1200 -50 1215
rect 2400 2385 2450 2400
rect 2400 1215 2410 2385
rect 2435 1215 2450 2385
rect 2400 1200 2450 1215
<< nsubdiff >>
rect -100 3695 -50 3710
rect -100 2525 -85 3695
rect -60 2525 -50 3695
rect -100 2510 -50 2525
rect 2400 3695 2450 3710
rect 2400 2525 2410 3695
rect 2435 2525 2450 3695
rect 2400 2510 2450 2525
<< psubdiffcont >>
rect -85 1215 -60 2385
rect 2410 1215 2435 2385
<< nsubdiffcont >>
rect -85 2525 -60 3695
rect 2410 2525 2435 3695
<< poly >>
rect -45 3755 100 3760
rect -45 3735 -35 3755
rect -15 3735 100 3755
rect -45 3730 100 3735
rect 0 3710 100 3730
rect 150 3755 2200 3760
rect 150 3735 415 3755
rect 435 3735 1915 3755
rect 1935 3735 2200 3755
rect 150 3725 2200 3735
rect 150 3710 250 3725
rect 300 3710 400 3725
rect 530 3710 630 3725
rect 660 3710 760 3725
rect 790 3710 890 3725
rect 920 3710 1020 3725
rect 1050 3710 1150 3725
rect 1200 3710 1300 3725
rect 1330 3710 1430 3725
rect 1460 3710 1560 3725
rect 1590 3710 1690 3725
rect 1720 3710 1820 3725
rect 1950 3710 2050 3725
rect 2100 3710 2200 3725
rect 2250 3755 2395 3760
rect 2250 3735 2365 3755
rect 2385 3735 2395 3755
rect 2250 3725 2395 3735
rect 2250 3710 2350 3725
rect 0 2495 100 2510
rect 150 2495 250 2510
rect 300 2495 400 2510
rect 530 2495 630 2510
rect 660 2495 760 2510
rect 790 2495 890 2510
rect 920 2495 1020 2510
rect 1050 2495 1150 2510
rect 1200 2495 1300 2510
rect 1330 2495 1430 2510
rect 1460 2495 1560 2510
rect 1590 2495 1690 2510
rect 1720 2495 1820 2510
rect 1950 2495 2050 2510
rect 2100 2495 2200 2510
rect 2250 2495 2350 2510
rect 300 2465 2050 2470
rect 300 2445 565 2465
rect 585 2445 865 2465
rect 885 2445 1465 2465
rect 1485 2445 1765 2465
rect 1785 2445 2050 2465
rect -45 2440 100 2445
rect -45 2420 -35 2440
rect -15 2420 100 2440
rect -45 2415 100 2420
rect 300 2440 2050 2445
rect 0 2400 100 2415
rect 150 2400 250 2415
rect 300 2400 400 2440
rect 450 2400 550 2440
rect 600 2400 700 2440
rect 750 2400 850 2440
rect 900 2400 1000 2440
rect 1050 2400 1150 2415
rect 1200 2400 1300 2415
rect 1350 2400 1450 2440
rect 1500 2400 1600 2440
rect 1650 2400 1750 2440
rect 1800 2400 1900 2440
rect 1950 2400 2050 2440
rect 2250 2440 2395 2445
rect 2250 2420 2365 2440
rect 2385 2420 2395 2440
rect 2250 2415 2395 2420
rect 2100 2400 2200 2415
rect 2250 2400 2350 2415
rect 0 1185 100 1200
rect 150 1180 250 1200
rect 300 1185 400 1200
rect 450 1185 550 1200
rect 600 1185 700 1200
rect 750 1185 850 1200
rect 900 1185 1000 1200
rect 1050 1185 1150 1200
rect 1200 1185 1300 1200
rect 1350 1185 1450 1200
rect 1500 1185 1600 1200
rect 1650 1185 1750 1200
rect 1800 1185 1900 1200
rect 1950 1185 2050 1200
rect 150 1160 160 1180
rect 240 1160 250 1180
rect 150 1155 250 1160
rect 1050 1180 1300 1185
rect 1050 1160 1165 1180
rect 1185 1160 1300 1180
rect 1050 1155 1300 1160
rect 2100 1180 2200 1200
rect 2250 1185 2350 1200
rect 2100 1160 2110 1180
rect 2190 1160 2200 1180
rect 2100 1155 2200 1160
<< polycont >>
rect -35 3735 -15 3755
rect 415 3735 435 3755
rect 1915 3735 1935 3755
rect 2365 3735 2385 3755
rect 565 2445 585 2465
rect 865 2445 885 2465
rect 1465 2445 1485 2465
rect 1765 2445 1785 2465
rect -35 2420 -15 2440
rect 2365 2420 2385 2440
rect 160 1160 240 1180
rect 1165 1160 1185 1180
rect 2110 1160 2190 1180
<< locali >>
rect -45 3755 -5 3760
rect -45 3735 -35 3755
rect -15 3735 -5 3755
rect -45 3705 -5 3735
rect 405 3755 445 3760
rect 405 3735 415 3755
rect 435 3735 445 3755
rect -95 3695 -5 3705
rect -95 2525 -85 3695
rect -60 2525 -40 3695
rect -15 2525 -5 3695
rect -95 2515 -5 2525
rect 105 3695 145 3705
rect 105 2525 115 3695
rect 135 2525 145 3695
rect 105 2495 145 2525
rect 255 3695 295 3705
rect 255 2525 265 3695
rect 285 2525 295 3695
rect 255 2515 295 2525
rect 405 3695 445 3735
rect 1905 3755 1945 3760
rect 1905 3735 1915 3755
rect 1935 3735 1945 3755
rect 405 2525 415 3695
rect 435 2525 445 3695
rect -100 2490 145 2495
rect -100 2470 105 2490
rect 135 2470 145 2490
rect -100 2465 145 2470
rect -45 2440 -5 2445
rect -45 2420 -35 2440
rect -15 2420 -5 2440
rect 405 2435 445 2525
rect 485 3695 525 3705
rect 485 2525 495 3695
rect 515 2525 525 3695
rect 485 2470 525 2525
rect 1155 3695 1195 3705
rect 1155 2525 1165 3695
rect 1185 2525 1195 3695
rect 1155 2515 1195 2525
rect 1825 3695 1865 3705
rect 1825 2525 1835 3695
rect 1855 2525 1865 3695
rect 1825 2470 1865 2525
rect 485 2465 595 2470
rect 485 2445 565 2465
rect 585 2445 595 2465
rect 485 2440 595 2445
rect -45 2395 -5 2420
rect -95 2385 -5 2395
rect -95 1215 -85 2385
rect -60 1215 -40 2385
rect -15 1215 -5 2385
rect -95 1205 -5 1215
rect 105 2415 445 2435
rect 105 2385 145 2415
rect 105 1215 115 2385
rect 135 1215 145 2385
rect 105 1205 145 1215
rect 255 2385 295 2395
rect 255 1215 265 2385
rect 285 1215 295 2385
rect 255 1205 295 1215
rect 405 2385 445 2395
rect 405 1215 415 2385
rect 435 1215 445 2385
rect 405 1185 445 1215
rect 555 2385 595 2440
rect 855 2465 895 2470
rect 855 2445 865 2465
rect 885 2445 895 2465
rect 555 1215 565 2385
rect 585 1215 595 2385
rect 555 1205 595 1215
rect 705 2385 745 2395
rect 705 1215 715 2385
rect 735 1215 745 2385
rect 705 1185 745 1215
rect 855 2385 895 2445
rect 1455 2465 1495 2470
rect 1455 2445 1465 2465
rect 1485 2445 1495 2465
rect 855 1215 865 2385
rect 885 1215 895 2385
rect 855 1205 895 1215
rect 1005 2385 1045 2395
rect 1005 1215 1015 2385
rect 1035 1215 1045 2385
rect 1005 1190 1045 1215
rect 1005 1185 1015 1190
rect 150 1180 250 1185
rect 150 1160 160 1180
rect 240 1160 250 1180
rect 405 1170 1015 1185
rect 1035 1170 1045 1190
rect 405 1165 1045 1170
rect 1155 2385 1195 2395
rect 1155 1215 1165 2385
rect 1185 1215 1195 2385
rect 1155 1180 1195 1215
rect 150 1155 250 1160
rect 1155 1160 1165 1180
rect 1185 1160 1195 1180
rect 1305 2385 1345 2395
rect 1305 1215 1315 2385
rect 1335 1215 1345 2385
rect 1305 1190 1345 1215
rect 1455 2385 1495 2445
rect 1755 2465 1865 2470
rect 1755 2445 1765 2465
rect 1785 2445 1865 2465
rect 1755 2440 1865 2445
rect 1905 3695 1945 3735
rect 2355 3755 2395 3760
rect 2355 3735 2365 3755
rect 2385 3735 2395 3755
rect 2355 3705 2395 3735
rect 1905 2525 1915 3695
rect 1935 2525 1945 3695
rect 1455 1215 1465 2385
rect 1485 1215 1495 2385
rect 1455 1205 1495 1215
rect 1605 2385 1645 2395
rect 1605 1215 1615 2385
rect 1635 1215 1645 2385
rect 1305 1170 1315 1190
rect 1335 1185 1345 1190
rect 1605 1185 1645 1215
rect 1755 2385 1795 2440
rect 1905 2435 1945 2525
rect 2055 3695 2095 3705
rect 2055 2525 2065 3695
rect 2085 2525 2095 3695
rect 2055 2515 2095 2525
rect 2205 3695 2245 3705
rect 2205 2525 2215 3695
rect 2235 2525 2245 3695
rect 2205 2515 2245 2525
rect 2355 3695 2445 3705
rect 2355 2525 2365 3695
rect 2390 2525 2410 3695
rect 2435 2525 2445 3695
rect 2355 2515 2445 2525
rect 2355 2440 2395 2445
rect 1905 2415 2245 2435
rect 1755 1215 1765 2385
rect 1785 1215 1795 2385
rect 1755 1205 1795 1215
rect 1905 2385 1945 2395
rect 1905 1215 1915 2385
rect 1935 1215 1945 2385
rect 1905 1185 1945 1215
rect 2055 2385 2095 2395
rect 2055 1215 2065 2385
rect 2085 1215 2095 2385
rect 2055 1205 2095 1215
rect 2205 2385 2245 2415
rect 2205 1215 2215 2385
rect 2235 1215 2245 2385
rect 2205 1205 2245 1215
rect 2355 2420 2365 2440
rect 2385 2420 2395 2440
rect 2355 2395 2395 2420
rect 2355 2385 2445 2395
rect 2355 1215 2365 2385
rect 2390 1215 2410 2385
rect 2435 1215 2445 2385
rect 2355 1205 2445 1215
rect 1335 1170 1945 1185
rect 1305 1165 1945 1170
rect 2100 1180 2200 1185
rect 1155 1155 1195 1160
rect 2100 1160 2110 1180
rect 2190 1160 2200 1180
rect 2100 1155 2200 1160
<< viali >>
rect -85 2525 -60 3695
rect -40 2525 -15 3695
rect 265 2525 285 3695
rect 105 2470 135 2490
rect 1165 2525 1185 3695
rect -85 1215 -60 2385
rect -40 1215 -15 2385
rect 265 1215 285 2385
rect 160 1160 240 1180
rect 1015 1170 1035 1190
rect 1165 2285 1185 2385
rect 1315 1170 1335 1190
rect 2065 2525 2085 3695
rect 2215 2525 2235 2625
rect 2365 2525 2390 3695
rect 2410 2525 2435 3695
rect 2065 1215 2085 2385
rect 2365 1215 2390 2385
rect 2410 1215 2435 2385
rect 2110 1160 2190 1180
<< metal1 >>
rect -95 3700 -5 3710
rect -95 2520 -90 3700
rect -60 2520 -40 3700
rect -10 2520 -5 3700
rect -95 2515 -5 2520
rect 255 3700 295 3705
rect 255 2520 260 3700
rect 290 2520 295 3700
rect 255 2515 295 2520
rect 1155 3700 1195 3705
rect 1155 2520 1160 3700
rect 1190 2520 1195 3700
rect 1155 2515 1195 2520
rect 2055 3700 2095 3705
rect 2055 2520 2060 3700
rect 2090 2520 2095 3700
rect 2355 3700 2445 3705
rect 2055 2515 2095 2520
rect 2205 2625 2245 2635
rect 2205 2525 2215 2625
rect 2235 2525 2245 2625
rect 2205 2495 2245 2525
rect 2355 2520 2360 3700
rect 2390 2520 2410 3700
rect 2440 2520 2445 3700
rect 2355 2515 2445 2520
rect 95 2490 2245 2495
rect 95 2470 105 2490
rect 135 2470 2245 2490
rect 95 2465 2245 2470
rect -95 2390 -5 2395
rect -95 1210 -90 2390
rect -55 1210 -40 2390
rect -10 1210 -5 2390
rect -95 1205 -5 1210
rect 255 2390 295 2395
rect 255 1210 260 2390
rect 290 1210 295 2390
rect 1155 2385 1195 2465
rect 1155 2285 1165 2385
rect 1185 2285 1195 2385
rect 1155 2275 1195 2285
rect 2055 2390 2095 2395
rect 255 1205 295 1210
rect 705 1215 1645 1245
rect 705 1185 745 1215
rect -100 1180 745 1185
rect -100 1160 160 1180
rect 240 1160 745 1180
rect 1005 1190 1345 1195
rect 1005 1170 1015 1190
rect 1035 1170 1315 1190
rect 1335 1170 1345 1190
rect 1005 1165 1345 1170
rect 1605 1185 1645 1215
rect 2055 1210 2060 2390
rect 2090 1210 2095 2390
rect 2055 1205 2095 1210
rect 2355 2390 2445 2395
rect 2355 1210 2360 2390
rect 2390 1210 2410 2390
rect 2440 1210 2445 2390
rect 2355 1205 2445 1210
rect 1605 1180 2200 1185
rect -100 1155 745 1160
rect 1605 1160 2110 1180
rect 2190 1160 2200 1180
rect 1605 1155 2200 1160
<< via1 >>
rect -90 3695 -60 3700
rect -90 2525 -85 3695
rect -85 2525 -60 3695
rect -90 2520 -60 2525
rect -40 3695 -10 3700
rect -40 2525 -15 3695
rect -15 2525 -10 3695
rect -40 2520 -10 2525
rect 260 3695 290 3700
rect 260 2525 265 3695
rect 265 2525 285 3695
rect 285 2525 290 3695
rect 260 2520 290 2525
rect 1160 3695 1190 3700
rect 1160 2525 1165 3695
rect 1165 2525 1185 3695
rect 1185 2525 1190 3695
rect 1160 2520 1190 2525
rect 2060 3695 2090 3700
rect 2060 2525 2065 3695
rect 2065 2525 2085 3695
rect 2085 2525 2090 3695
rect 2060 2520 2090 2525
rect 2360 3695 2390 3700
rect 2360 2525 2365 3695
rect 2365 2525 2390 3695
rect 2360 2520 2390 2525
rect 2410 3695 2440 3700
rect 2410 2525 2435 3695
rect 2435 2525 2440 3695
rect 2410 2520 2440 2525
rect -90 2385 -55 2390
rect -90 1215 -85 2385
rect -85 1215 -60 2385
rect -60 1215 -55 2385
rect -90 1210 -55 1215
rect -40 2385 -10 2390
rect -40 1215 -15 2385
rect -15 1215 -10 2385
rect -40 1210 -10 1215
rect 260 2385 290 2390
rect 260 1215 265 2385
rect 265 1215 285 2385
rect 285 1215 290 2385
rect 260 1210 290 1215
rect 2060 2385 2090 2390
rect 2060 1215 2065 2385
rect 2065 1215 2085 2385
rect 2085 1215 2090 2385
rect 2060 1210 2090 1215
rect 2360 2385 2390 2390
rect 2360 1215 2365 2385
rect 2365 1215 2390 2385
rect 2360 1210 2390 1215
rect 2410 2385 2440 2390
rect 2410 1215 2435 2385
rect 2435 1215 2440 2385
rect 2410 1210 2440 1215
<< metal2 >>
rect -95 3705 -5 3710
rect -100 3700 2450 3705
rect -100 2520 -90 3700
rect -60 2520 -40 3700
rect -10 2520 260 3700
rect 290 2520 1160 3700
rect 1190 2520 2060 3700
rect 2090 2520 2360 3700
rect 2390 2520 2410 3700
rect 2440 2520 2450 3700
rect -100 2515 2450 2520
rect -100 2390 2450 2395
rect -100 1210 -90 2390
rect -55 1210 -40 2390
rect -10 1210 260 2390
rect 290 1210 2060 2390
rect 2090 1210 2360 2390
rect 2390 1210 2410 2390
rect 2440 1210 2450 2390
rect -100 1205 2450 1210
<< labels >>
rlabel metal1 -100 1170 -100 1170 7 Vbn
port 1 w
rlabel metal2 -100 1800 -100 1800 7 VN
port 2 w
rlabel locali -100 2480 -100 2480 7 Vgate
port 3 w
rlabel metal2 -100 3110 -100 3110 7 VP
port 4 w
<< end >>
