magic
tech sky130A
timestamp 1699571337
<< error_p >>
rect 2905 0 2955 1200
rect 3055 0 3105 1200
rect 3205 0 3255 1200
rect 3355 0 3405 1200
rect 3505 0 3555 1200
rect 3655 0 3705 1200
<< nmos >>
rect -155 0 -55 1200
rect -5 0 95 1200
rect 145 0 245 1200
rect 295 0 395 1200
rect 445 0 545 1200
rect 675 0 775 1200
rect 825 0 925 1200
rect 975 0 1075 1200
rect 1125 0 1225 1200
rect 1455 0 1555 1200
rect 1605 0 1705 1200
rect 1755 0 1855 1200
rect 1905 0 2005 1200
rect 2055 0 2155 1200
rect 2205 0 2305 1200
rect 2355 0 2455 1200
rect 2505 0 2605 1200
rect 2655 0 2755 1200
rect 2805 0 2905 1200
rect 2955 0 3055 1200
rect 3105 0 3205 1200
rect 3255 0 3355 1200
rect 3405 0 3505 1200
rect 3555 0 3655 1200
rect 3705 0 3805 1200
rect 3855 0 3955 1200
rect 4005 0 4105 1200
rect 4155 0 4255 1200
rect 4305 0 4405 1200
rect 4455 0 4555 1200
rect 4605 0 4705 1200
rect 4755 0 4855 1200
rect 4905 0 5005 1200
rect 5055 0 5155 1200
<< ndiff >>
rect -205 1185 -155 1200
rect -205 15 -190 1185
rect -170 15 -155 1185
rect -205 0 -155 15
rect -55 1185 -5 1200
rect -55 15 -40 1185
rect -20 15 -5 1185
rect -55 0 -5 15
rect 95 1185 145 1200
rect 95 15 110 1185
rect 130 15 145 1185
rect 95 0 145 15
rect 245 1185 295 1200
rect 245 15 260 1185
rect 280 15 295 1185
rect 245 0 295 15
rect 395 1185 445 1200
rect 395 15 410 1185
rect 430 15 445 1185
rect 395 0 445 15
rect 545 1185 595 1200
rect 545 15 560 1185
rect 580 15 595 1185
rect 545 0 595 15
rect 625 1185 675 1200
rect 625 15 640 1185
rect 660 15 675 1185
rect 625 0 675 15
rect 775 1185 825 1200
rect 775 15 790 1185
rect 810 15 825 1185
rect 775 0 825 15
rect 925 1185 975 1200
rect 925 15 940 1185
rect 960 15 975 1185
rect 925 0 975 15
rect 1075 1185 1125 1200
rect 1075 15 1090 1185
rect 1110 15 1125 1185
rect 1075 0 1125 15
rect 1225 1185 1275 1200
rect 1225 15 1240 1185
rect 1260 15 1275 1185
rect 1225 0 1275 15
rect 1405 1185 1455 1200
rect 1405 15 1420 1185
rect 1440 15 1455 1185
rect 1405 0 1455 15
rect 1555 1185 1605 1200
rect 1555 15 1570 1185
rect 1590 15 1605 1185
rect 1555 0 1605 15
rect 1705 1185 1755 1200
rect 1705 15 1720 1185
rect 1740 15 1755 1185
rect 1705 0 1755 15
rect 1855 1185 1905 1200
rect 1855 15 1870 1185
rect 1890 15 1905 1185
rect 1855 0 1905 15
rect 2005 1185 2055 1200
rect 2005 15 2020 1185
rect 2040 15 2055 1185
rect 2005 0 2055 15
rect 2155 1185 2205 1200
rect 2155 15 2170 1185
rect 2190 15 2205 1185
rect 2155 0 2205 15
rect 2305 1185 2355 1200
rect 2305 15 2320 1185
rect 2340 15 2355 1185
rect 2305 0 2355 15
rect 2455 1185 2505 1200
rect 2455 15 2470 1185
rect 2490 15 2505 1185
rect 2455 0 2505 15
rect 2605 1185 2655 1200
rect 2605 15 2620 1185
rect 2640 15 2655 1185
rect 2605 0 2655 15
rect 2755 1185 2805 1200
rect 2755 15 2770 1185
rect 2790 15 2805 1185
rect 2755 0 2805 15
rect 2905 1185 2955 1200
rect 2905 15 2920 1185
rect 2940 15 2955 1185
rect 2905 0 2955 15
rect 3055 1185 3105 1200
rect 3055 15 3070 1185
rect 3090 15 3105 1185
rect 3055 0 3105 15
rect 3205 1185 3255 1200
rect 3205 15 3220 1185
rect 3240 15 3255 1185
rect 3205 0 3255 15
rect 3355 1185 3405 1200
rect 3355 15 3370 1185
rect 3390 15 3405 1185
rect 3355 0 3405 15
rect 3505 1185 3555 1200
rect 3505 15 3520 1185
rect 3540 15 3555 1185
rect 3505 0 3555 15
rect 3655 1185 3705 1200
rect 3655 15 3670 1185
rect 3690 15 3705 1185
rect 3655 0 3705 15
rect 3805 1185 3855 1200
rect 3805 15 3820 1185
rect 3840 15 3855 1185
rect 3805 0 3855 15
rect 3955 1185 4005 1200
rect 3955 15 3970 1185
rect 3990 15 4005 1185
rect 3955 0 4005 15
rect 4105 1185 4155 1200
rect 4105 15 4120 1185
rect 4140 15 4155 1185
rect 4105 0 4155 15
rect 4255 1185 4305 1200
rect 4255 15 4270 1185
rect 4290 15 4305 1185
rect 4255 0 4305 15
rect 4405 1185 4455 1200
rect 4405 15 4420 1185
rect 4440 15 4455 1185
rect 4405 0 4455 15
rect 4555 1185 4605 1200
rect 4555 15 4570 1185
rect 4590 15 4605 1185
rect 4555 0 4605 15
rect 4705 1185 4755 1200
rect 4705 15 4720 1185
rect 4740 15 4755 1185
rect 4705 0 4755 15
rect 4855 1185 4905 1200
rect 4855 15 4870 1185
rect 4890 15 4905 1185
rect 4855 0 4905 15
rect 5005 1185 5055 1200
rect 5005 15 5020 1185
rect 5040 15 5055 1185
rect 5005 0 5055 15
rect 5155 1185 5205 1200
rect 5155 15 5170 1185
rect 5190 15 5205 1185
rect 5155 0 5205 15
<< ndiffc >>
rect -190 15 -170 1185
rect -40 15 -20 1185
rect 110 15 130 1185
rect 260 15 280 1185
rect 410 15 430 1185
rect 560 15 580 1185
rect 640 15 660 1185
rect 790 15 810 1185
rect 940 15 960 1185
rect 1090 15 1110 1185
rect 1240 15 1260 1185
rect 1420 15 1440 1185
rect 1570 15 1590 1185
rect 1720 15 1740 1185
rect 1870 15 1890 1185
rect 2020 15 2040 1185
rect 2170 15 2190 1185
rect 2320 15 2340 1185
rect 2470 15 2490 1185
rect 2620 15 2640 1185
rect 2770 15 2790 1185
rect 2920 15 2940 1185
rect 3070 15 3090 1185
rect 3220 15 3240 1185
rect 3370 15 3390 1185
rect 3520 15 3540 1185
rect 3670 15 3690 1185
rect 3820 15 3840 1185
rect 3970 15 3990 1185
rect 4120 15 4140 1185
rect 4270 15 4290 1185
rect 4420 15 4440 1185
rect 4570 15 4590 1185
rect 4720 15 4740 1185
rect 4870 15 4890 1185
rect 5020 15 5040 1185
rect 5170 15 5190 1185
<< psubdiff >>
rect -255 1185 -205 1200
rect -255 15 -240 1185
rect -220 15 -205 1185
rect -255 0 -205 15
rect 1355 1185 1405 1200
rect 1355 15 1370 1185
rect 1390 15 1405 1185
rect 1355 0 1405 15
rect 5205 1185 5255 1200
rect 5205 15 5220 1185
rect 5240 15 5255 1185
rect 5205 0 5255 15
<< psubdiffcont >>
rect -240 15 -220 1185
rect 1370 15 1390 1185
rect 5220 15 5240 1185
<< poly >>
rect 680 1240 720 1250
rect 680 1225 690 1240
rect 675 1220 690 1225
rect 710 1230 720 1240
rect 2610 1245 2650 1255
rect 2610 1235 2620 1245
rect 710 1220 1225 1230
rect 675 1215 1225 1220
rect 1605 1215 2455 1230
rect -155 1200 -55 1215
rect -5 1200 95 1215
rect 145 1200 245 1215
rect 295 1200 395 1215
rect 445 1200 545 1215
rect 675 1200 775 1215
rect 825 1200 925 1215
rect 975 1200 1075 1215
rect 1125 1200 1225 1215
rect 1455 1200 1555 1215
rect 1605 1200 1705 1215
rect 1755 1200 1855 1215
rect 1905 1200 2005 1215
rect 2055 1200 2155 1215
rect 2205 1200 2305 1215
rect 2355 1200 2455 1215
rect 2505 1225 2620 1235
rect 2640 1235 2650 1245
rect 2910 1245 2950 1255
rect 2910 1235 2920 1245
rect 2640 1225 2920 1235
rect 2940 1235 2950 1245
rect 3040 1240 3420 1255
rect 3040 1235 3055 1240
rect 2940 1225 3055 1235
rect 2505 1215 3055 1225
rect 3405 1235 3420 1240
rect 3510 1245 3550 1255
rect 3510 1235 3520 1245
rect 3405 1225 3520 1235
rect 3540 1235 3550 1245
rect 3810 1245 3850 1255
rect 3810 1235 3820 1245
rect 3540 1225 3820 1235
rect 3840 1235 3850 1245
rect 3840 1225 3955 1235
rect 3405 1215 3955 1225
rect 2505 1200 2605 1215
rect 2655 1200 2755 1215
rect 2805 1200 2905 1215
rect 2955 1200 3055 1215
rect 3105 1200 3205 1215
rect 3255 1200 3355 1215
rect 3405 1200 3505 1215
rect 3555 1200 3655 1215
rect 3705 1200 3805 1215
rect 3855 1200 3955 1215
rect 4005 1200 4105 1215
rect 4155 1200 4255 1215
rect 4305 1200 4405 1215
rect 4455 1200 4555 1215
rect 4605 1200 4705 1215
rect 4755 1200 4855 1215
rect 4905 1200 5005 1215
rect 5055 1200 5155 1215
rect -155 -15 -55 0
rect -5 -10 95 0
rect 145 -10 245 0
rect 295 -10 395 0
rect 445 -10 545 0
rect -5 -20 545 -10
rect 675 -15 775 0
rect 825 -15 925 0
rect 975 -15 1075 0
rect 1125 -15 1225 0
rect 1455 -15 1555 0
rect 1605 -15 1705 0
rect 1755 -15 1855 0
rect 1905 -15 2005 0
rect 2055 -15 2155 0
rect 2205 -15 2305 0
rect 2355 -15 2455 0
rect -5 -25 260 -20
rect 250 -40 260 -25
rect 280 -25 545 -20
rect 1455 -20 1495 -15
rect 280 -40 290 -25
rect 1455 -40 1465 -20
rect 1485 -40 1495 -20
rect 250 -50 290 -40
rect 870 -50 1030 -40
rect 1455 -50 1495 -40
rect 1755 -20 1795 -15
rect 1755 -40 1765 -20
rect 1785 -40 1795 -20
rect 1755 -50 1795 -40
rect 1965 -20 2005 -15
rect 1965 -40 1975 -20
rect 1995 -40 2005 -20
rect 2505 -30 2605 0
rect 2655 -15 2755 0
rect 2805 -15 2905 0
rect 2655 -30 2905 -15
rect 2955 -30 3055 0
rect 3105 -15 3205 0
rect 3255 -15 3355 0
rect 3405 -30 3505 0
rect 3555 -15 3655 0
rect 3705 -15 3805 0
rect 3555 -30 3805 -15
rect 3855 -30 3955 0
rect 4005 -15 4105 0
rect 4155 -15 4255 0
rect 4305 -15 4405 0
rect 4455 -15 4555 0
rect 4605 -15 4705 0
rect 4755 -15 4855 0
rect 4905 -15 5005 0
rect 5055 -15 5155 0
rect 1965 -50 2005 -40
rect 250 -110 265 -50
rect 870 -70 880 -50
rect 900 -55 1000 -50
rect 900 -70 910 -55
rect 870 -80 910 -70
rect 990 -70 1000 -55
rect 1020 -70 1030 -50
rect 990 -80 1030 -70
rect 250 -120 290 -110
rect 250 -140 260 -120
rect 280 -140 290 -120
rect 250 -150 290 -140
<< polycont >>
rect 690 1220 710 1240
rect 2620 1225 2640 1245
rect 2920 1225 2940 1245
rect 3520 1225 3540 1245
rect 3820 1225 3840 1245
rect 260 -40 280 -20
rect 1465 -40 1485 -20
rect 1765 -40 1785 -20
rect 1975 -40 1995 -20
rect 880 -70 900 -50
rect 1000 -70 1020 -50
rect 260 -140 280 -120
<< locali >>
rect 680 1240 720 1250
rect 550 1220 690 1240
rect 710 1220 720 1240
rect 550 1215 720 1220
rect -250 1185 -160 1195
rect -250 15 -240 1185
rect -220 15 -190 1185
rect -170 15 -160 1185
rect -250 5 -160 15
rect -50 1185 -10 1195
rect -50 15 -40 1185
rect -20 15 -10 1185
rect -50 -70 -10 15
rect 100 1185 140 1195
rect 100 15 110 1185
rect 130 15 140 1185
rect 100 5 140 15
rect 250 1185 290 1195
rect 250 15 260 1185
rect 280 15 290 1185
rect 250 -20 290 15
rect 400 1185 440 1195
rect 400 15 410 1185
rect 430 15 440 1185
rect 400 5 440 15
rect 550 1185 590 1215
rect 680 1210 720 1215
rect 2610 1245 2650 1255
rect 2610 1225 2620 1245
rect 2640 1225 2650 1245
rect 550 15 560 1185
rect 580 15 590 1185
rect 250 -40 260 -20
rect 280 -40 290 -20
rect 250 -50 290 -40
rect 550 -70 590 15
rect 630 1185 670 1195
rect 630 15 640 1185
rect 660 15 670 1185
rect 630 -40 670 15
rect 780 1185 820 1195
rect 780 15 790 1185
rect 810 15 820 1185
rect 780 5 820 15
rect 930 1185 970 1195
rect 930 15 940 1185
rect 960 15 970 1185
rect 630 -50 910 -40
rect 630 -60 880 -50
rect -50 -90 590 -70
rect 870 -70 880 -60
rect 900 -70 910 -50
rect 870 -80 910 -70
rect 250 -120 290 -110
rect 250 -140 260 -120
rect 280 -140 290 -120
rect 930 -140 970 15
rect 1080 1185 1120 1195
rect 1080 15 1090 1185
rect 1110 15 1120 1185
rect 1080 5 1120 15
rect 1230 1185 1270 1195
rect 1230 15 1240 1185
rect 1260 15 1270 1185
rect 1230 -40 1270 15
rect 1360 1185 1450 1195
rect 1360 15 1370 1185
rect 1390 15 1420 1185
rect 1440 15 1450 1185
rect 1360 5 1450 15
rect 1560 1185 1600 1195
rect 1560 15 1570 1185
rect 1590 15 1600 1185
rect 1560 5 1600 15
rect 1710 1185 1750 1195
rect 1710 15 1720 1185
rect 1740 15 1750 1185
rect 990 -50 1270 -40
rect 1410 -10 1450 5
rect 1710 -10 1750 15
rect 1860 1185 1900 1195
rect 1860 15 1870 1185
rect 1890 15 1900 1185
rect 1860 5 1900 15
rect 2010 1185 2050 1195
rect 2010 15 2020 1185
rect 2040 15 2050 1185
rect 2010 -10 2050 15
rect 2160 1185 2200 1195
rect 2160 15 2170 1185
rect 2190 15 2200 1185
rect 2160 5 2200 15
rect 2310 1185 2350 1195
rect 2310 15 2320 1185
rect 2340 15 2350 1185
rect 2310 5 2350 15
rect 2460 1185 2500 1195
rect 2460 15 2470 1185
rect 2490 15 2500 1185
rect 1410 -20 1495 -10
rect 1410 -40 1465 -20
rect 1485 -40 1495 -20
rect 1410 -50 1495 -40
rect 1710 -20 1795 -10
rect 1710 -40 1765 -20
rect 1785 -40 1795 -20
rect 1710 -50 1795 -40
rect 1965 -20 2050 -10
rect 1965 -40 1975 -20
rect 1995 -40 2050 -20
rect 1965 -50 2050 -40
rect 2460 -30 2500 15
rect 2610 1185 2650 1225
rect 2910 1245 2950 1255
rect 2910 1225 2920 1245
rect 2940 1225 2950 1245
rect 2610 15 2620 1185
rect 2640 15 2650 1185
rect 2610 5 2650 15
rect 2760 1185 2800 1195
rect 2760 15 2770 1185
rect 2790 15 2800 1185
rect 2760 -30 2800 15
rect 2910 1185 2950 1225
rect 3510 1245 3550 1255
rect 3510 1225 3520 1245
rect 3540 1225 3550 1245
rect 2910 15 2920 1185
rect 2940 15 2950 1185
rect 2910 5 2950 15
rect 3060 1185 3100 1195
rect 3060 15 3070 1185
rect 3090 15 3100 1185
rect 3060 -30 3100 15
rect 3210 1185 3250 1195
rect 3210 15 3220 1185
rect 3240 15 3250 1185
rect 3210 5 3250 15
rect 3360 1185 3400 1195
rect 3360 15 3370 1185
rect 3390 15 3400 1185
rect 3360 -30 3400 15
rect 3510 1185 3550 1225
rect 3810 1245 3850 1255
rect 3810 1225 3820 1245
rect 3840 1225 3850 1245
rect 3510 15 3520 1185
rect 3540 15 3550 1185
rect 3510 5 3550 15
rect 3660 1185 3700 1195
rect 3660 15 3670 1185
rect 3690 15 3700 1185
rect 3660 -30 3700 15
rect 3810 1185 3850 1225
rect 3810 15 3820 1185
rect 3840 15 3850 1185
rect 3810 5 3850 15
rect 3960 1185 4000 1195
rect 3960 15 3970 1185
rect 3990 15 4000 1185
rect 3960 -30 4000 15
rect 4110 1185 4150 1195
rect 4110 15 4120 1185
rect 4140 15 4150 1185
rect 4110 5 4150 15
rect 4260 1185 4300 1195
rect 4260 15 4270 1185
rect 4290 15 4300 1185
rect 4260 5 4300 15
rect 4410 1185 4450 1195
rect 4410 15 4420 1185
rect 4440 15 4450 1185
rect 4410 5 4450 15
rect 4560 1185 4600 1195
rect 4560 15 4570 1185
rect 4590 15 4600 1185
rect 4560 5 4600 15
rect 4710 1185 4750 1195
rect 4710 15 4720 1185
rect 4740 15 4750 1185
rect 4710 5 4750 15
rect 4860 1185 4900 1195
rect 4860 15 4870 1185
rect 4890 15 4900 1185
rect 4860 5 4900 15
rect 5010 1185 5050 1195
rect 5010 15 5020 1185
rect 5040 15 5050 1185
rect 5010 5 5050 15
rect 5160 1185 5250 1195
rect 5160 15 5170 1185
rect 5190 15 5220 1185
rect 5240 15 5250 1185
rect 5160 5 5250 15
rect 2460 -50 4000 -30
rect 990 -70 1000 -50
rect 1020 -60 1270 -50
rect 1020 -70 1030 -60
rect 990 -80 1030 -70
rect 250 -150 290 -140
<< end >>
