magic
tech sky130A
timestamp 1699634882
<< poly >>
rect 10874 1353 11196 1360
rect 10874 1335 11166 1353
rect 11186 1335 11196 1353
rect 10874 1330 11196 1335
<< polycont >>
rect 11166 1335 11186 1353
<< locali >>
rect 5730 2337 5805 2370
rect 5730 1460 5755 2337
rect 5647 1439 5755 1460
rect 11152 1353 11191 1360
rect 11152 1335 11166 1353
rect 11186 1335 11191 1353
rect 11152 1330 11191 1335
use big  big_0
timestamp 1699632857
transform 1 0 275 0 1 1565
box -275 -1545 5375 1255
use cascode_biasgen  cascode_biasgen_0
timestamp 1699590019
transform 1 0 11291 0 1 -1135
box -120 1155 2470 3760
use dac  dac_0
timestamp 1699634024
transform 0 1 8241 -1 0 2630
box -101 -2457 2602 2659
<< end >>
