magic
tech sky130A
timestamp 1699659720
<< nwell >>
rect 11170 2525 11175 2530
rect 5540 2185 5565 2345
rect 5570 2185 5580 2345
rect 11115 2250 11175 2525
rect 5515 2095 5590 2185
rect 5540 2070 5565 2095
rect 5570 2070 5580 2095
rect 5535 1540 5585 1740
rect 11115 1670 11175 1945
rect 11170 1665 11175 1670
rect 5755 1020 5805 1160
rect 11110 755 11160 895
rect 5735 560 5785 580
rect 5715 460 5785 560
rect 5735 440 5785 460
<< nsubdiff >>
rect 5735 1125 5785 1140
rect 5735 1055 5750 1125
rect 5770 1055 5785 1125
rect 5735 1040 5785 1055
rect 11090 860 11140 875
rect 11090 790 11105 860
rect 11125 790 11140 860
rect 11090 775 11140 790
rect 5715 545 5765 560
rect 5715 475 5730 545
rect 5750 475 5765 545
rect 5715 460 5765 475
<< nsubdiffcont >>
rect 5750 1055 5770 1125
rect 11105 790 11125 860
rect 5730 475 5750 545
<< poly >>
rect 10920 1950 10960 1960
rect 10920 1930 10930 1950
rect 10950 1930 10960 1950
rect 10920 1920 10960 1930
rect 10920 1880 10935 1920
rect 5775 1860 5830 1870
rect 10855 1865 10935 1880
rect 5775 1840 5785 1860
rect 5805 1840 5830 1860
rect 5775 1830 5830 1840
rect 5775 1660 5830 1670
rect 5775 1640 5785 1660
rect 5805 1640 5830 1660
rect 5775 1630 5830 1640
rect 10855 1630 10915 1645
rect 10900 1570 10915 1630
rect 10900 1560 10940 1570
rect 10900 1540 10910 1560
rect 10930 1540 10940 1560
rect 10900 1530 10940 1540
rect 10874 1353 11196 1360
rect 10874 1335 11166 1353
rect 11186 1335 11196 1353
rect 10874 1330 11196 1335
rect 5775 660 5830 670
rect 5775 640 5785 660
rect 5805 640 5830 660
rect 5775 630 5830 640
rect 10855 610 10895 620
rect 10855 590 10865 610
rect 10885 590 10895 610
rect 10855 580 10895 590
rect 5785 460 5830 470
rect 5785 440 5795 460
rect 5815 440 5830 460
rect 5785 430 5830 440
<< polycont >>
rect 10930 1930 10950 1950
rect 5785 1840 5805 1860
rect 5785 1640 5805 1660
rect 10910 1540 10930 1560
rect 11166 1335 11186 1353
rect 5785 640 5805 660
rect 10865 590 10885 610
rect 5795 440 5815 460
<< locali >>
rect 5545 2340 5785 2370
rect 5545 1440 5565 2340
rect 10920 2230 11025 2250
rect 5690 2050 5795 2070
rect 5775 1870 5795 2050
rect 10920 1960 10940 2230
rect 10920 1950 10960 1960
rect 10920 1930 10930 1950
rect 10950 1930 10960 1950
rect 10920 1920 10960 1930
rect 5775 1860 5815 1870
rect 5775 1840 5785 1860
rect 5805 1840 5815 1860
rect 5775 1830 5815 1840
rect 5775 1660 5815 1670
rect 5775 1640 5785 1660
rect 5805 1640 5815 1660
rect 5775 1630 5815 1640
rect 10920 1650 11030 1670
rect 5775 1465 5795 1630
rect 10920 1570 10940 1650
rect 10900 1560 10940 1570
rect 10900 1540 10910 1560
rect 10930 1540 10940 1560
rect 10900 1530 10940 1540
rect 5690 1445 5795 1465
rect 11152 1353 11191 1360
rect 11152 1335 11166 1353
rect 11186 1335 11191 1353
rect 11152 1330 11191 1335
rect 5690 1125 5780 1135
rect 5690 1055 5750 1125
rect 5770 1055 5780 1125
rect 5690 1045 5780 1055
rect 5625 865 5795 885
rect 5775 670 5795 865
rect 11045 860 11135 870
rect 11045 790 11105 860
rect 11125 790 11135 860
rect 11045 780 11135 790
rect 5775 660 5815 670
rect 5775 640 5785 660
rect 5805 640 5815 660
rect 5775 630 5815 640
rect 10855 610 10985 620
rect 10855 590 10865 610
rect 10885 600 10985 610
rect 10885 590 10895 600
rect 10855 580 10895 590
rect 5710 545 5760 555
rect 5710 475 5730 545
rect 5750 475 5760 545
rect 5710 465 5760 475
rect 5785 460 5825 470
rect 5785 440 5795 460
rect 5815 440 5825 460
rect 5785 430 5825 440
rect 5785 305 5805 430
rect 5635 285 5805 305
<< viali >>
rect 5750 1055 5770 1125
rect 11105 790 11125 860
rect 5730 475 5750 545
<< metal1 >>
rect 5525 2485 11090 2500
rect 5525 2425 5540 2485
rect 5760 2425 11090 2485
rect 5525 2410 11090 2425
rect 10865 2275 10960 2365
rect 5505 2095 5590 2185
rect 5505 1580 5545 2095
rect 10865 2030 10900 2275
rect 5715 1940 10900 2030
rect 10865 1785 10900 1940
rect 10865 1695 10965 1785
rect 5505 1490 5595 1580
rect 5505 1000 5545 1490
rect 5690 1130 5780 1135
rect 5690 1050 5745 1130
rect 5775 1050 5780 1130
rect 5690 1045 5780 1050
rect 5505 910 5590 1000
rect 5505 420 5545 910
rect 10865 735 10900 1695
rect 11045 865 11150 870
rect 11045 785 11100 865
rect 11130 785 11150 865
rect 11045 780 11150 785
rect 10865 645 10940 735
rect 5710 550 5760 555
rect 5710 470 5725 550
rect 5755 470 5760 550
rect 5710 465 5760 470
rect 5505 330 5590 420
rect 10865 50 10900 645
rect 11110 295 11150 780
rect 11110 100 11115 295
rect 11145 100 11150 295
rect 11110 95 11150 100
rect 10865 20 11200 50
<< via1 >>
rect 5540 2425 5760 2485
rect 5745 1125 5775 1130
rect 5745 1055 5750 1125
rect 5750 1055 5770 1125
rect 5770 1055 5775 1125
rect 5745 1050 5775 1055
rect 11100 860 11130 865
rect 11100 790 11105 860
rect 11105 790 11125 860
rect 11125 790 11130 860
rect 11100 785 11130 790
rect 5725 545 5755 550
rect 5725 475 5730 545
rect 5730 475 5750 545
rect 5750 475 5755 545
rect 5725 470 5755 475
rect 11115 100 11145 295
<< metal2 >>
rect 5525 2485 5780 2500
rect 5525 2425 5540 2485
rect 5760 2425 5780 2485
rect 5525 2410 5780 2425
rect 11090 2410 11200 2500
rect 5520 2230 5755 2320
rect 5585 1805 5845 2185
rect 10840 1985 11130 2365
rect 11090 1830 11200 1920
rect 5525 1625 5755 1715
rect 5430 1135 5520 1570
rect 5585 1200 5845 1580
rect 10840 1405 11130 1785
rect 11190 1385 11200 1390
rect 11230 1385 11240 1390
rect 11190 1360 11240 1385
rect 11045 1320 11240 1360
rect 5430 1130 5780 1135
rect 5430 1050 5745 1130
rect 5775 1050 5780 1130
rect 5430 1045 5780 1050
rect 5430 555 5520 1045
rect 5560 620 5845 1000
rect 11045 870 11085 1320
rect 11045 865 11135 870
rect 11045 785 11100 865
rect 11130 785 11135 865
rect 11045 780 11135 785
rect 5430 550 5760 555
rect 5430 470 5725 550
rect 5755 470 5760 550
rect 5430 465 5760 470
rect 5235 60 5845 420
rect 10840 355 11195 735
rect 10840 295 11150 300
rect 10840 100 11115 295
rect 11145 100 11150 295
rect 10840 95 11150 100
use big  big_0
timestamp 1699632857
transform 1 0 170 0 1 1565
box -275 -1545 5375 1255
use cascode_biasgen  cascode_biasgen_0
timestamp 1699636225
transform 1 0 11291 0 1 -1135
box -120 1155 2470 3760
use dac  dac_0
timestamp 1699653726
transform 0 1 8241 -1 0 2630
box -101 -2457 2602 2659
use mux_tall  mux_tall_0
timestamp 1699649434
transform 1 0 10860 0 1 2130
box 75 -165 295 395
use mux_tall  mux_tall_1
timestamp 1699649434
transform 1 0 10860 0 1 1550
box 75 -165 295 395
use mux_tall  mux_tall_2
timestamp 1699649434
transform 1 0 10815 0 1 500
box 75 -165 295 395
use mux_tall  mux_tall_3
timestamp 1699649434
transform 1 0 5440 0 1 185
box 75 -165 295 395
use mux_tall  mux_tall_4
timestamp 1699649434
transform 1 0 5460 0 1 765
box 75 -165 295 395
use mux_tall  mux_tall_5
timestamp 1699649434
transform 1 0 5485 0 1 1345
box 75 -165 295 395
use mux_tall  mux_tall_6
timestamp 1699649434
transform 1 0 5485 0 1 1950
box 75 -165 295 395
<< end >>
