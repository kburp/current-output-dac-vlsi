magic
tech sky130A
timestamp 1699632857
<< nwell >>
rect -275 -25 5375 1235
<< nmos >>
rect -155 -1510 -55 -310
rect -5 -1510 95 -310
rect 225 -1510 325 -310
rect 375 -1510 475 -310
rect 525 -1510 625 -310
rect 675 -1510 775 -310
rect 825 -1510 925 -310
rect 975 -1510 1075 -310
rect 1125 -1510 1225 -310
rect 1275 -1510 1375 -310
rect 1425 -1510 1525 -310
rect 1575 -1510 1675 -310
rect 1725 -1510 1825 -310
rect 1875 -1510 1975 -310
rect 2025 -1510 2125 -310
rect 2175 -1510 2275 -310
rect 2325 -1510 2425 -310
rect 2475 -1510 2575 -310
rect 2755 -1510 2855 -310
rect 2985 -1510 3085 -310
rect 3135 -1510 3235 -310
rect 3285 -1510 3385 -310
rect 3435 -1510 3535 -310
rect 3665 -1510 3765 -310
rect 3815 -1510 3915 -310
rect 3965 -1510 4065 -310
rect 4115 -1510 4215 -310
rect 4265 -1510 4365 -310
rect 4415 -1510 4515 -310
rect 4565 -1510 4665 -310
rect 4715 -1510 4815 -310
rect 4865 -1510 4965 -310
<< pmos >>
rect -155 0 -55 1200
rect -5 0 95 1200
rect 145 0 245 1200
rect 295 0 395 1200
rect 445 0 545 1200
rect 675 0 775 1200
rect 825 0 925 1200
rect 975 0 1075 1200
rect 1125 0 1225 1200
rect 1355 0 1455 1200
rect 1505 0 1605 1200
rect 1655 0 1755 1200
rect 1805 0 1905 1200
rect 1955 0 2055 1200
rect 2105 0 2205 1200
rect 2355 0 2455 1200
rect 2505 0 2605 1200
rect 2655 0 2755 1200
rect 2805 0 2905 1200
rect 2955 0 3055 1200
rect 3105 0 3205 1200
rect 3255 0 3355 1200
rect 3405 0 3505 1200
rect 3555 0 3655 1200
rect 3705 0 3805 1200
rect 3855 0 3955 1200
rect 4005 0 4105 1200
rect 4255 0 4355 1200
rect 4405 0 4505 1200
rect 4555 0 4655 1200
rect 4705 0 4805 1200
rect 4855 0 4955 1200
rect 5005 0 5105 1200
rect 5155 0 5255 1200
<< ndiff >>
rect -205 -325 -155 -310
rect -205 -1495 -190 -325
rect -170 -1495 -155 -325
rect -205 -1510 -155 -1495
rect -55 -325 -5 -310
rect -55 -1495 -40 -325
rect -20 -1495 -5 -325
rect -55 -1510 -5 -1495
rect 95 -325 145 -310
rect 95 -1495 110 -325
rect 130 -1495 145 -325
rect 95 -1510 145 -1495
rect 175 -325 225 -310
rect 175 -1495 190 -325
rect 210 -1495 225 -325
rect 175 -1510 225 -1495
rect 325 -325 375 -310
rect 325 -1495 340 -325
rect 360 -1495 375 -325
rect 325 -1510 375 -1495
rect 475 -325 525 -310
rect 475 -1495 490 -325
rect 510 -1495 525 -325
rect 475 -1510 525 -1495
rect 625 -325 675 -310
rect 625 -1495 640 -325
rect 660 -1495 675 -325
rect 625 -1510 675 -1495
rect 775 -325 825 -310
rect 775 -1495 790 -325
rect 810 -1495 825 -325
rect 775 -1510 825 -1495
rect 925 -325 975 -310
rect 925 -1495 940 -325
rect 960 -1495 975 -325
rect 925 -1510 975 -1495
rect 1075 -325 1125 -310
rect 1075 -1495 1090 -325
rect 1110 -1495 1125 -325
rect 1075 -1510 1125 -1495
rect 1225 -325 1275 -310
rect 1225 -1495 1240 -325
rect 1260 -1495 1275 -325
rect 1225 -1510 1275 -1495
rect 1375 -325 1425 -310
rect 1375 -1495 1390 -325
rect 1410 -1495 1425 -325
rect 1375 -1510 1425 -1495
rect 1525 -325 1575 -310
rect 1525 -1495 1540 -325
rect 1560 -1495 1575 -325
rect 1525 -1510 1575 -1495
rect 1675 -325 1725 -310
rect 1675 -1495 1690 -325
rect 1710 -1495 1725 -325
rect 1675 -1510 1725 -1495
rect 1825 -325 1875 -310
rect 1825 -1495 1840 -325
rect 1860 -1495 1875 -325
rect 1825 -1510 1875 -1495
rect 1975 -325 2025 -310
rect 1975 -1495 1990 -325
rect 2010 -1495 2025 -325
rect 1975 -1510 2025 -1495
rect 2125 -325 2175 -310
rect 2125 -1495 2140 -325
rect 2160 -1495 2175 -325
rect 2125 -1510 2175 -1495
rect 2275 -325 2325 -310
rect 2275 -1495 2290 -325
rect 2310 -1495 2325 -325
rect 2275 -1510 2325 -1495
rect 2425 -325 2475 -310
rect 2425 -1495 2440 -325
rect 2460 -1495 2475 -325
rect 2425 -1510 2475 -1495
rect 2575 -325 2625 -310
rect 2575 -1495 2590 -325
rect 2610 -1495 2625 -325
rect 2575 -1510 2625 -1495
rect 2705 -325 2755 -310
rect 2705 -1495 2720 -325
rect 2740 -1495 2755 -325
rect 2705 -1510 2755 -1495
rect 2855 -325 2905 -310
rect 2855 -1495 2870 -325
rect 2890 -1495 2905 -325
rect 2855 -1510 2905 -1495
rect 2935 -325 2985 -310
rect 2935 -1495 2950 -325
rect 2970 -1495 2985 -325
rect 2935 -1510 2985 -1495
rect 3085 -325 3135 -310
rect 3085 -1495 3100 -325
rect 3120 -1495 3135 -325
rect 3085 -1510 3135 -1495
rect 3235 -325 3285 -310
rect 3235 -1495 3250 -325
rect 3270 -1495 3285 -325
rect 3235 -1510 3285 -1495
rect 3385 -325 3435 -310
rect 3385 -1495 3400 -325
rect 3420 -1495 3435 -325
rect 3385 -1510 3435 -1495
rect 3535 -325 3585 -310
rect 3535 -1495 3550 -325
rect 3570 -1495 3585 -325
rect 3535 -1510 3585 -1495
rect 3615 -325 3665 -310
rect 3615 -1495 3630 -325
rect 3650 -1495 3665 -325
rect 3615 -1510 3665 -1495
rect 3765 -325 3815 -310
rect 3765 -1495 3780 -325
rect 3800 -1495 3815 -325
rect 3765 -1510 3815 -1495
rect 3915 -325 3965 -310
rect 3915 -1495 3930 -325
rect 3950 -1495 3965 -325
rect 3915 -1510 3965 -1495
rect 4065 -325 4115 -310
rect 4065 -1495 4080 -325
rect 4100 -1495 4115 -325
rect 4065 -1510 4115 -1495
rect 4215 -325 4265 -310
rect 4215 -1495 4230 -325
rect 4250 -1495 4265 -325
rect 4215 -1510 4265 -1495
rect 4365 -325 4415 -310
rect 4365 -1495 4380 -325
rect 4400 -1495 4415 -325
rect 4365 -1510 4415 -1495
rect 4515 -325 4565 -310
rect 4515 -1495 4530 -325
rect 4550 -1495 4565 -325
rect 4515 -1510 4565 -1495
rect 4665 -325 4715 -310
rect 4665 -1495 4680 -325
rect 4700 -1495 4715 -325
rect 4665 -1510 4715 -1495
rect 4815 -325 4865 -310
rect 4815 -1495 4830 -325
rect 4850 -1495 4865 -325
rect 4815 -1510 4865 -1495
rect 4965 -325 5015 -310
rect 4965 -1495 4980 -325
rect 5000 -1495 5015 -325
rect 4965 -1510 5015 -1495
<< pdiff >>
rect -205 1185 -155 1200
rect -205 15 -190 1185
rect -170 15 -155 1185
rect -205 0 -155 15
rect -55 1185 -5 1200
rect -55 15 -40 1185
rect -20 15 -5 1185
rect -55 0 -5 15
rect 95 1185 145 1200
rect 95 15 110 1185
rect 130 15 145 1185
rect 95 0 145 15
rect 245 1185 295 1200
rect 245 15 260 1185
rect 280 15 295 1185
rect 245 0 295 15
rect 395 1185 445 1200
rect 395 15 410 1185
rect 430 15 445 1185
rect 395 0 445 15
rect 545 1185 595 1200
rect 545 15 560 1185
rect 580 15 595 1185
rect 545 0 595 15
rect 625 1185 675 1200
rect 625 15 640 1185
rect 660 15 675 1185
rect 625 0 675 15
rect 775 1185 825 1200
rect 775 15 790 1185
rect 810 15 825 1185
rect 775 0 825 15
rect 925 1185 975 1200
rect 925 15 940 1185
rect 960 15 975 1185
rect 925 0 975 15
rect 1075 1185 1125 1200
rect 1075 15 1090 1185
rect 1110 15 1125 1185
rect 1075 0 1125 15
rect 1225 1185 1275 1200
rect 1225 15 1240 1185
rect 1260 15 1275 1185
rect 1225 0 1275 15
rect 1305 1185 1355 1200
rect 1305 15 1320 1185
rect 1340 15 1355 1185
rect 1305 0 1355 15
rect 1455 1185 1505 1200
rect 1455 15 1470 1185
rect 1490 15 1505 1185
rect 1455 0 1505 15
rect 1605 1185 1655 1200
rect 1605 15 1620 1185
rect 1640 15 1655 1185
rect 1605 0 1655 15
rect 1755 1185 1805 1200
rect 1755 15 1770 1185
rect 1790 15 1805 1185
rect 1755 0 1805 15
rect 1905 1185 1955 1200
rect 1905 15 1920 1185
rect 1940 15 1955 1185
rect 1905 0 1955 15
rect 2055 1185 2105 1200
rect 2055 15 2070 1185
rect 2090 15 2105 1185
rect 2055 0 2105 15
rect 2205 1185 2255 1200
rect 2305 1185 2355 1200
rect 2205 15 2220 1185
rect 2240 15 2255 1185
rect 2305 15 2320 1185
rect 2340 15 2355 1185
rect 2205 0 2255 15
rect 2305 0 2355 15
rect 2455 1185 2505 1200
rect 2455 15 2470 1185
rect 2490 15 2505 1185
rect 2455 0 2505 15
rect 2605 1185 2655 1200
rect 2605 15 2620 1185
rect 2640 15 2655 1185
rect 2605 0 2655 15
rect 2755 1185 2805 1200
rect 2755 15 2770 1185
rect 2790 15 2805 1185
rect 2755 0 2805 15
rect 2905 1185 2955 1200
rect 2905 15 2920 1185
rect 2940 15 2955 1185
rect 2905 0 2955 15
rect 3055 1185 3105 1200
rect 3055 15 3070 1185
rect 3090 15 3105 1185
rect 3055 0 3105 15
rect 3205 1185 3255 1200
rect 3205 15 3220 1185
rect 3240 15 3255 1185
rect 3205 0 3255 15
rect 3355 1185 3405 1200
rect 3355 15 3370 1185
rect 3390 15 3405 1185
rect 3355 0 3405 15
rect 3505 1185 3555 1200
rect 3505 15 3520 1185
rect 3540 15 3555 1185
rect 3505 0 3555 15
rect 3655 1185 3705 1200
rect 3655 15 3670 1185
rect 3690 15 3705 1185
rect 3655 0 3705 15
rect 3805 1185 3855 1200
rect 3805 15 3820 1185
rect 3840 15 3855 1185
rect 3805 0 3855 15
rect 3955 1185 4005 1200
rect 3955 15 3970 1185
rect 3990 15 4005 1185
rect 3955 0 4005 15
rect 4105 1185 4155 1200
rect 4205 1185 4255 1200
rect 4105 15 4120 1185
rect 4140 15 4155 1185
rect 4205 15 4220 1185
rect 4240 15 4255 1185
rect 4105 0 4155 15
rect 4205 0 4255 15
rect 4355 1185 4405 1200
rect 4355 15 4370 1185
rect 4390 15 4405 1185
rect 4355 0 4405 15
rect 4505 1185 4555 1200
rect 4505 15 4520 1185
rect 4540 15 4555 1185
rect 4505 0 4555 15
rect 4655 1185 4705 1200
rect 4655 15 4670 1185
rect 4690 15 4705 1185
rect 4655 0 4705 15
rect 4805 1185 4855 1200
rect 4805 15 4820 1185
rect 4840 15 4855 1185
rect 4805 0 4855 15
rect 4955 1185 5005 1200
rect 4955 15 4970 1185
rect 4990 15 5005 1185
rect 4955 0 5005 15
rect 5105 1185 5155 1200
rect 5105 15 5120 1185
rect 5140 15 5155 1185
rect 5105 0 5155 15
rect 5255 1185 5305 1200
rect 5255 15 5270 1185
rect 5290 15 5305 1185
rect 5255 0 5305 15
<< ndiffc >>
rect -190 -1495 -170 -325
rect -40 -1495 -20 -325
rect 110 -1495 130 -325
rect 190 -1495 210 -325
rect 340 -1495 360 -325
rect 490 -1495 510 -325
rect 640 -1495 660 -325
rect 790 -1495 810 -325
rect 940 -1495 960 -325
rect 1090 -1495 1110 -325
rect 1240 -1495 1260 -325
rect 1390 -1495 1410 -325
rect 1540 -1495 1560 -325
rect 1690 -1495 1710 -325
rect 1840 -1495 1860 -325
rect 1990 -1495 2010 -325
rect 2140 -1495 2160 -325
rect 2290 -1495 2310 -325
rect 2440 -1495 2460 -325
rect 2590 -1495 2610 -325
rect 2720 -1495 2740 -325
rect 2870 -1495 2890 -325
rect 2950 -1495 2970 -325
rect 3100 -1495 3120 -325
rect 3250 -1495 3270 -325
rect 3400 -1495 3420 -325
rect 3550 -1495 3570 -325
rect 3630 -1495 3650 -325
rect 3780 -1495 3800 -325
rect 3930 -1495 3950 -325
rect 4080 -1495 4100 -325
rect 4230 -1495 4250 -325
rect 4380 -1495 4400 -325
rect 4530 -1495 4550 -325
rect 4680 -1495 4700 -325
rect 4830 -1495 4850 -325
rect 4980 -1495 5000 -325
<< pdiffc >>
rect -190 15 -170 1185
rect -40 15 -20 1185
rect 110 15 130 1185
rect 260 15 280 1185
rect 410 15 430 1185
rect 560 15 580 1185
rect 640 15 660 1185
rect 790 15 810 1185
rect 940 15 960 1185
rect 1090 15 1110 1185
rect 1240 15 1260 1185
rect 1320 15 1340 1185
rect 1470 15 1490 1185
rect 1620 15 1640 1185
rect 1770 15 1790 1185
rect 1920 15 1940 1185
rect 2070 15 2090 1185
rect 2220 15 2240 1185
rect 2320 15 2340 1185
rect 2470 15 2490 1185
rect 2620 15 2640 1185
rect 2770 15 2790 1185
rect 2920 15 2940 1185
rect 3070 15 3090 1185
rect 3220 15 3240 1185
rect 3370 15 3390 1185
rect 3520 15 3540 1185
rect 3670 15 3690 1185
rect 3820 15 3840 1185
rect 3970 15 3990 1185
rect 4120 15 4140 1185
rect 4220 15 4240 1185
rect 4370 15 4390 1185
rect 4520 15 4540 1185
rect 4670 15 4690 1185
rect 4820 15 4840 1185
rect 4970 15 4990 1185
rect 5120 15 5140 1185
rect 5270 15 5290 1185
<< psubdiff >>
rect -255 -325 -205 -310
rect -255 -1495 -240 -325
rect -220 -1495 -205 -325
rect -255 -1510 -205 -1495
rect 2655 -325 2705 -310
rect 2655 -1495 2670 -325
rect 2690 -1495 2705 -325
rect 2655 -1510 2705 -1495
rect 5015 -325 5065 -310
rect 5015 -1495 5030 -325
rect 5050 -1495 5065 -325
rect 5015 -1510 5065 -1495
<< nsubdiff >>
rect -255 1185 -205 1200
rect -255 15 -240 1185
rect -220 15 -205 1185
rect -255 0 -205 15
rect 2255 1185 2305 1200
rect 2255 15 2270 1185
rect 2290 15 2305 1185
rect 2255 0 2305 15
rect 4155 1185 4205 1200
rect 4155 15 4170 1185
rect 4190 15 4205 1185
rect 4155 0 4205 15
rect 5305 1185 5355 1200
rect 5305 15 5320 1185
rect 5340 15 5355 1185
rect 5305 0 5355 15
<< psubdiffcont >>
rect -240 -1495 -220 -325
rect 2670 -1495 2690 -325
rect 5030 -1495 5050 -325
<< nsubdiffcont >>
rect -240 15 -220 1185
rect 2270 15 2290 1185
rect 4170 15 4190 1185
rect 5320 15 5340 1185
<< poly >>
rect 675 1245 715 1255
rect 675 1225 685 1245
rect 705 1230 715 1245
rect 1655 1245 1695 1255
rect 1655 1230 1665 1245
rect 705 1225 1225 1230
rect 675 1215 1225 1225
rect 1505 1225 1665 1230
rect 1685 1230 1695 1245
rect 1865 1245 1905 1255
rect 1865 1230 1875 1245
rect 1685 1225 1875 1230
rect 1895 1230 1905 1245
rect 2610 1245 2650 1255
rect 2610 1230 2620 1245
rect 1895 1225 2455 1230
rect 1505 1215 2455 1225
rect -155 1200 -55 1215
rect -5 1200 95 1215
rect 145 1200 245 1215
rect 295 1200 395 1215
rect 445 1200 545 1215
rect 675 1200 775 1215
rect 825 1200 925 1215
rect 975 1200 1075 1215
rect 1125 1200 1225 1215
rect 1355 1200 1455 1215
rect 1505 1200 1605 1215
rect 1655 1200 1755 1215
rect 1805 1200 1905 1215
rect 1955 1200 2055 1215
rect 2105 1200 2205 1215
rect 2355 1200 2455 1215
rect 2505 1225 2620 1230
rect 2640 1230 2650 1245
rect 2910 1245 2950 1255
rect 2910 1230 2920 1245
rect 2640 1225 2920 1230
rect 2940 1230 2950 1245
rect 3040 1240 3420 1255
rect 3040 1230 3055 1240
rect 2940 1225 3055 1230
rect 2505 1215 3055 1225
rect 3405 1230 3420 1240
rect 3510 1245 3550 1255
rect 3510 1230 3520 1245
rect 3405 1225 3520 1230
rect 3540 1230 3550 1245
rect 3810 1245 3850 1255
rect 3810 1230 3820 1245
rect 3540 1225 3820 1230
rect 3840 1230 3850 1245
rect 4555 1245 4595 1255
rect 4555 1230 4565 1245
rect 3840 1225 3955 1230
rect 3405 1215 3955 1225
rect 2505 1200 2605 1215
rect 2655 1200 2755 1215
rect 2805 1200 2905 1215
rect 2955 1200 3055 1215
rect 3105 1200 3205 1215
rect 3255 1200 3355 1215
rect 3405 1200 3505 1215
rect 3555 1200 3655 1215
rect 3705 1200 3805 1215
rect 3855 1200 3955 1215
rect 4005 1225 4565 1230
rect 4585 1230 4595 1245
rect 4765 1245 4805 1255
rect 4765 1230 4775 1245
rect 4585 1225 4775 1230
rect 4795 1230 4805 1245
rect 4795 1225 4955 1230
rect 4005 1215 4955 1225
rect 4005 1200 4105 1215
rect 4255 1200 4355 1215
rect 4405 1200 4505 1215
rect 4555 1200 4655 1215
rect 4705 1200 4805 1215
rect 4855 1200 4955 1215
rect 5005 1200 5105 1215
rect 5155 1200 5255 1215
rect -155 -15 -55 0
rect -5 -10 95 0
rect 145 -10 245 0
rect 295 -10 395 0
rect 445 -10 545 0
rect -155 -25 -115 -15
rect -5 -25 545 -10
rect 675 -15 775 0
rect 825 -15 925 0
rect 975 -15 1075 0
rect 1125 -15 1225 0
rect 1355 -15 1455 0
rect 1505 -15 1605 0
rect 1655 -15 1755 0
rect 1805 -15 1905 0
rect 1955 -15 2055 0
rect 2105 -15 2205 0
rect 2355 -15 2455 0
rect 2505 -15 2605 0
rect 2655 -15 2755 0
rect 2805 -15 2905 0
rect 2955 -15 3055 0
rect 3105 -15 3205 0
rect 1355 -25 1395 -15
rect -155 -45 -145 -25
rect -125 -45 -115 -25
rect -155 -55 -115 -45
rect 250 -45 260 -25
rect 280 -45 290 -25
rect 250 -55 290 -45
rect 1355 -45 1365 -25
rect 1385 -45 1395 -25
rect 1355 -55 1395 -45
rect 2400 -25 2440 -15
rect 2400 -45 2410 -25
rect 2430 -45 2440 -25
rect 2400 -55 2440 -45
rect 250 -115 265 -55
rect 250 -125 290 -115
rect 250 -145 260 -125
rect 280 -145 290 -125
rect 250 -155 290 -145
rect 570 -140 610 -130
rect 570 -160 580 -140
rect 600 -155 610 -140
rect 690 -140 730 -130
rect 3190 -135 3205 -15
rect 690 -155 700 -140
rect 600 -160 700 -155
rect 720 -160 730 -140
rect 570 -170 730 -160
rect 3165 -145 3205 -135
rect 3165 -165 3175 -145
rect 3195 -165 3205 -145
rect 3165 -175 3205 -165
rect 3255 -15 3355 0
rect 3405 -15 3505 0
rect 3555 -15 3655 0
rect 3705 -15 3805 0
rect 3855 -15 3955 0
rect 4005 -15 4105 0
rect 4255 -15 4355 0
rect 4405 -15 4505 0
rect 4555 -15 4655 0
rect 4705 -15 4805 0
rect 4855 -15 4955 0
rect 5005 -15 5105 0
rect 5155 -15 5255 0
rect 3255 -135 3270 -15
rect 3255 -145 3295 -135
rect 3255 -165 3265 -145
rect 3285 -165 3295 -145
rect 3255 -175 3295 -165
rect 3640 -175 3655 -15
rect 4020 -25 4060 -15
rect 4020 -45 4030 -25
rect 4050 -45 4060 -25
rect 5065 -25 5105 -15
rect 4020 -55 4060 -45
rect 4450 -50 4610 -40
rect 4450 -70 4460 -50
rect 4480 -55 4580 -50
rect 4480 -70 4490 -55
rect 4450 -80 4490 -70
rect 4570 -70 4580 -55
rect 4600 -70 4610 -50
rect 5065 -45 5075 -25
rect 5095 -45 5105 -25
rect 5065 -55 5105 -45
rect 5215 -25 5255 -15
rect 5215 -45 5225 -25
rect 5245 -45 5255 -25
rect 5215 -55 5255 -45
rect 4570 -80 4610 -70
rect 4450 -115 4610 -105
rect 4450 -135 4460 -115
rect 4480 -120 4580 -115
rect 4480 -135 4490 -120
rect 4450 -145 4490 -135
rect 4570 -135 4580 -120
rect 4600 -135 4610 -115
rect 4570 -145 4610 -135
rect 3620 -185 3660 -175
rect 570 -205 730 -195
rect 570 -225 580 -205
rect 600 -210 700 -205
rect 600 -225 610 -210
rect 570 -235 610 -225
rect 690 -225 700 -210
rect 720 -225 730 -205
rect 3620 -205 3630 -185
rect 3650 -205 3660 -185
rect 3620 -215 3660 -205
rect 690 -235 730 -225
rect -155 -265 -115 -255
rect -155 -285 -145 -265
rect -125 -285 -115 -265
rect 330 -265 370 -255
rect 330 -280 340 -265
rect -155 -295 -115 -285
rect -5 -285 340 -280
rect 360 -280 370 -265
rect 630 -265 670 -255
rect 630 -280 640 -265
rect 360 -285 640 -280
rect 660 -280 670 -265
rect 930 -265 970 -255
rect 930 -280 940 -265
rect 660 -285 940 -280
rect 960 -280 970 -265
rect 1230 -265 1270 -255
rect 1230 -280 1240 -265
rect 960 -285 1240 -280
rect 1260 -280 1270 -265
rect 1530 -265 1570 -255
rect 1530 -280 1540 -265
rect 1260 -285 1540 -280
rect 1560 -280 1570 -265
rect 1830 -265 1870 -255
rect 1830 -280 1840 -265
rect 1560 -285 1840 -280
rect 1860 -280 1870 -265
rect 2130 -265 2170 -255
rect 2130 -280 2140 -265
rect 1860 -285 2140 -280
rect 2160 -280 2170 -265
rect 2430 -265 2470 -255
rect 2430 -280 2440 -265
rect 2160 -285 2440 -280
rect 2460 -280 2470 -265
rect 3240 -265 3280 -255
rect 3240 -280 3250 -265
rect 2460 -285 2855 -280
rect -5 -295 2855 -285
rect -155 -310 -55 -295
rect -5 -310 95 -295
rect 225 -310 325 -295
rect 375 -310 475 -295
rect 525 -310 625 -295
rect 675 -310 775 -295
rect 825 -310 925 -295
rect 975 -310 1075 -295
rect 1125 -310 1225 -295
rect 1275 -310 1375 -295
rect 1425 -310 1525 -295
rect 1575 -310 1675 -295
rect 1725 -310 1825 -295
rect 1875 -310 1975 -295
rect 2025 -310 2125 -295
rect 2175 -310 2275 -295
rect 2325 -310 2425 -295
rect 2475 -310 2575 -295
rect 2755 -310 2855 -295
rect 2985 -285 3250 -280
rect 3270 -280 3280 -265
rect 3680 -265 3720 -255
rect 3680 -280 3690 -265
rect 3270 -285 3535 -280
rect 2985 -295 3535 -285
rect 2985 -310 3085 -295
rect 3135 -310 3235 -295
rect 3285 -310 3385 -295
rect 3435 -310 3535 -295
rect 3665 -285 3690 -280
rect 3710 -280 3720 -265
rect 4925 -265 4965 -255
rect 3710 -285 4815 -280
rect 3665 -295 4815 -285
rect 4925 -285 4935 -265
rect 4955 -285 4965 -265
rect 4925 -295 4965 -285
rect 3665 -310 3765 -295
rect 3815 -310 3915 -295
rect 3965 -310 4065 -295
rect 4115 -310 4215 -295
rect 4265 -310 4365 -295
rect 4415 -310 4515 -295
rect 4565 -310 4665 -295
rect 4715 -310 4815 -295
rect 4865 -310 4965 -295
rect -155 -1525 -55 -1510
rect -5 -1525 95 -1510
rect 225 -1525 325 -1510
rect 375 -1525 475 -1510
rect 525 -1525 625 -1510
rect 675 -1525 775 -1510
rect 825 -1525 925 -1510
rect 975 -1525 1075 -1510
rect 1125 -1525 1225 -1510
rect 1275 -1525 1375 -1510
rect 1425 -1525 1525 -1510
rect 1575 -1525 1675 -1510
rect 1725 -1525 1825 -1510
rect 1875 -1525 1975 -1510
rect 2025 -1525 2125 -1510
rect 2175 -1525 2275 -1510
rect 2325 -1525 2425 -1510
rect 2475 -1525 2575 -1510
rect 2755 -1525 2855 -1510
rect 2985 -1525 3085 -1510
rect 3135 -1525 3235 -1510
rect 3285 -1525 3385 -1510
rect 3435 -1525 3535 -1510
rect 3665 -1525 3765 -1510
rect 3815 -1525 3915 -1510
rect 3965 -1525 4065 -1510
rect 4115 -1525 4215 -1510
rect 4265 -1525 4365 -1510
rect 4415 -1525 4515 -1510
rect 4565 -1525 4665 -1510
rect 4715 -1525 4815 -1510
rect 4865 -1525 4965 -1510
<< polycont >>
rect 685 1225 705 1245
rect 1665 1225 1685 1245
rect 1875 1225 1895 1245
rect 2620 1225 2640 1245
rect 2920 1225 2940 1245
rect 3520 1225 3540 1245
rect 3820 1225 3840 1245
rect 4565 1225 4585 1245
rect 4775 1225 4795 1245
rect -145 -45 -125 -25
rect 260 -45 280 -25
rect 1365 -45 1385 -25
rect 2410 -45 2430 -25
rect 260 -145 280 -125
rect 580 -160 600 -140
rect 700 -160 720 -140
rect 3175 -165 3195 -145
rect 3265 -165 3285 -145
rect 4030 -45 4050 -25
rect 4460 -70 4480 -50
rect 4580 -70 4600 -50
rect 5075 -45 5095 -25
rect 5225 -45 5245 -25
rect 4460 -135 4480 -115
rect 4580 -135 4600 -115
rect 580 -225 600 -205
rect 700 -225 720 -205
rect 3630 -205 3650 -185
rect -145 -285 -125 -265
rect 340 -285 360 -265
rect 640 -285 660 -265
rect 940 -285 960 -265
rect 1240 -285 1260 -265
rect 1540 -285 1560 -265
rect 1840 -285 1860 -265
rect 2140 -285 2160 -265
rect 2440 -285 2460 -265
rect 3250 -285 3270 -265
rect 3690 -285 3710 -265
rect 4935 -285 4955 -265
<< locali >>
rect 675 1245 715 1255
rect 675 1240 685 1245
rect 550 1225 685 1240
rect 705 1225 715 1245
rect 550 1215 715 1225
rect 1610 1245 1695 1255
rect 1610 1225 1665 1245
rect 1685 1225 1695 1245
rect 1610 1215 1695 1225
rect 1865 1245 1950 1255
rect 1865 1225 1875 1245
rect 1895 1225 1950 1245
rect 1865 1215 1950 1225
rect -250 1185 -160 1195
rect -250 15 -240 1185
rect -220 15 -190 1185
rect -170 15 -160 1185
rect -250 5 -160 15
rect -200 -15 -160 5
rect -50 1185 -10 1195
rect -50 15 -40 1185
rect -20 15 -10 1185
rect -200 -25 -115 -15
rect -200 -45 -145 -25
rect -125 -45 -115 -25
rect -200 -55 -115 -45
rect -50 -75 -10 15
rect 100 1185 140 1195
rect 100 15 110 1185
rect 130 15 140 1185
rect 100 5 140 15
rect 250 1185 290 1195
rect 250 15 260 1185
rect 280 15 290 1185
rect 250 -25 290 15
rect 400 1185 440 1195
rect 400 15 410 1185
rect 430 15 440 1185
rect 400 5 440 15
rect 550 1185 590 1215
rect 550 15 560 1185
rect 580 15 590 1185
rect 250 -45 260 -25
rect 280 -45 290 -25
rect 250 -55 290 -45
rect 550 -75 590 15
rect -50 -95 590 -75
rect 250 -125 290 -115
rect 250 -145 260 -125
rect 280 -145 290 -125
rect 250 -155 290 -145
rect 570 -130 590 -95
rect 630 1185 670 1195
rect 630 15 640 1185
rect 660 15 670 1185
rect 630 -40 670 15
rect 780 1185 820 1195
rect 780 15 790 1185
rect 810 15 820 1185
rect 780 5 820 15
rect 930 1185 970 1195
rect 930 15 940 1185
rect 960 15 970 1185
rect 930 5 970 15
rect 1080 1185 1120 1195
rect 1080 15 1090 1185
rect 1110 15 1120 1185
rect 1080 5 1120 15
rect 1230 1185 1270 1195
rect 1230 15 1240 1185
rect 1260 15 1270 1185
rect 1230 -40 1270 15
rect 1305 1185 1350 1195
rect 1305 15 1320 1185
rect 1340 15 1350 1185
rect 1305 5 1350 15
rect 630 -60 1270 -40
rect 1310 -15 1350 5
rect 1460 1185 1500 1195
rect 1460 15 1470 1185
rect 1490 15 1500 1185
rect 1310 -25 1395 -15
rect 1310 -45 1365 -25
rect 1385 -45 1395 -25
rect 1310 -55 1395 -45
rect 570 -140 610 -130
rect 250 -215 270 -155
rect 570 -160 580 -140
rect 600 -160 610 -140
rect 570 -170 610 -160
rect 570 -205 610 -195
rect 570 -215 580 -205
rect -50 -225 580 -215
rect 600 -225 610 -205
rect -50 -235 610 -225
rect -200 -265 -115 -255
rect -200 -285 -145 -265
rect -125 -285 -115 -265
rect -200 -295 -115 -285
rect -200 -315 -160 -295
rect -50 -315 -10 -235
rect 330 -265 370 -255
rect 330 -285 340 -265
rect 360 -285 370 -265
rect -250 -325 -160 -315
rect -250 -1495 -240 -325
rect -220 -1495 -190 -325
rect -170 -1495 -160 -325
rect -250 -1505 -160 -1495
rect -55 -325 -10 -315
rect -55 -1495 -40 -325
rect -20 -1495 -10 -325
rect -55 -1505 -10 -1495
rect 100 -325 140 -315
rect 100 -1495 110 -325
rect 130 -1495 140 -325
rect 100 -1505 140 -1495
rect 180 -325 220 -315
rect 180 -1495 190 -325
rect 210 -1495 220 -325
rect 180 -1525 220 -1495
rect 330 -325 370 -285
rect 630 -265 670 -60
rect 1375 -95 1395 -55
rect 1460 -55 1500 15
rect 1610 1185 1650 1215
rect 1610 15 1620 1185
rect 1640 15 1650 1185
rect 1610 5 1650 15
rect 1760 1185 1800 1195
rect 1760 15 1770 1185
rect 1790 15 1800 1185
rect 1760 -55 1800 15
rect 1910 1185 1950 1215
rect 2610 1245 2650 1255
rect 2610 1225 2620 1245
rect 2640 1225 2650 1245
rect 1910 15 1920 1185
rect 1940 15 1950 1185
rect 1910 5 1950 15
rect 2060 1185 2100 1195
rect 2060 15 2070 1185
rect 2090 15 2100 1185
rect 2060 -55 2100 15
rect 2210 1185 2350 1195
rect 2210 15 2220 1185
rect 2240 15 2270 1185
rect 2290 15 2320 1185
rect 2340 15 2350 1185
rect 2210 5 2350 15
rect 2460 1185 2500 1195
rect 2460 15 2470 1185
rect 2490 15 2500 1185
rect 2460 -15 2500 15
rect 2610 1185 2650 1225
rect 2910 1245 2950 1255
rect 2910 1225 2920 1245
rect 2940 1225 2950 1245
rect 2610 15 2620 1185
rect 2640 15 2650 1185
rect 2610 5 2650 15
rect 2760 1185 2800 1195
rect 2760 15 2770 1185
rect 2790 15 2800 1185
rect 2760 -15 2800 15
rect 2910 1185 2950 1225
rect 2910 15 2920 1185
rect 2940 15 2950 1185
rect 2910 5 2950 15
rect 3060 1185 3100 1195
rect 3060 15 3070 1185
rect 3090 15 3100 1185
rect 3060 -15 3100 15
rect 3210 1185 3250 1255
rect 3510 1245 3550 1255
rect 3510 1225 3520 1245
rect 3540 1225 3550 1245
rect 3210 15 3220 1185
rect 3240 15 3250 1185
rect 3210 5 3250 15
rect 3360 1185 3400 1195
rect 3360 15 3370 1185
rect 3390 15 3400 1185
rect 3360 -15 3400 15
rect 3510 1185 3550 1225
rect 3810 1245 3850 1255
rect 3810 1225 3820 1245
rect 3840 1225 3850 1245
rect 3510 15 3520 1185
rect 3540 15 3550 1185
rect 3510 5 3550 15
rect 3660 1185 3700 1195
rect 3660 15 3670 1185
rect 3690 15 3700 1185
rect 3660 -15 3700 15
rect 3810 1185 3850 1225
rect 4510 1245 4595 1255
rect 4510 1225 4565 1245
rect 4585 1225 4595 1245
rect 4510 1215 4595 1225
rect 4765 1245 4850 1255
rect 4765 1225 4775 1245
rect 4795 1225 4850 1245
rect 4765 1215 4850 1225
rect 3810 15 3820 1185
rect 3840 15 3850 1185
rect 3810 5 3850 15
rect 3960 1185 4000 1195
rect 3960 15 3970 1185
rect 3990 15 4000 1185
rect 3960 -15 4000 15
rect 4110 1185 4250 1195
rect 4110 15 4120 1185
rect 4140 15 4170 1185
rect 4190 15 4220 1185
rect 4240 15 4250 1185
rect 4110 5 4250 15
rect 4360 1185 4400 1195
rect 4360 15 4370 1185
rect 4390 15 4400 1185
rect 2400 -25 2440 -15
rect 2400 -45 2410 -25
rect 2430 -45 2440 -25
rect 2460 -35 4000 -15
rect 4020 -25 4060 -15
rect 2400 -55 2440 -45
rect 4020 -45 4030 -25
rect 4050 -45 4060 -25
rect 4020 -55 4060 -45
rect 4360 -55 4400 15
rect 4510 1185 4550 1215
rect 4510 15 4520 1185
rect 4540 15 4550 1185
rect 4450 -50 4490 -40
rect 4450 -55 4460 -50
rect 1460 -75 2380 -55
rect 2420 -75 4040 -55
rect 4080 -70 4460 -55
rect 4480 -70 4490 -50
rect 4080 -75 4490 -70
rect 2360 -95 2380 -75
rect 4080 -95 4100 -75
rect 4450 -80 4490 -75
rect 1375 -115 2340 -95
rect 2360 -115 4100 -95
rect 4120 -115 4490 -105
rect 690 -140 730 -130
rect 690 -160 700 -140
rect 720 -150 730 -140
rect 2320 -135 2340 -115
rect 4120 -125 4460 -115
rect 4120 -135 4140 -125
rect 2320 -145 4140 -135
rect 4450 -135 4460 -125
rect 4480 -135 4490 -115
rect 4450 -145 4490 -135
rect 720 -160 770 -150
rect 2320 -155 3175 -145
rect 690 -170 770 -160
rect 750 -175 770 -170
rect 3165 -165 3175 -155
rect 3195 -155 3265 -145
rect 3195 -165 3205 -155
rect 3165 -175 3205 -165
rect 3255 -165 3265 -155
rect 3285 -155 4140 -145
rect 3285 -165 3295 -155
rect 3255 -175 3295 -165
rect 750 -195 2980 -175
rect 690 -205 730 -195
rect 690 -225 700 -205
rect 720 -215 730 -205
rect 2940 -215 2980 -195
rect 3620 -185 3660 -175
rect 3620 -205 3630 -185
rect 3650 -205 3660 -185
rect 720 -225 2900 -215
rect 690 -235 2900 -225
rect 630 -285 640 -265
rect 660 -285 670 -265
rect 330 -1495 340 -325
rect 360 -1495 370 -325
rect 330 -1505 370 -1495
rect 480 -325 520 -315
rect 480 -1495 490 -325
rect 510 -1495 520 -325
rect 480 -1525 520 -1495
rect 630 -325 670 -285
rect 930 -265 970 -255
rect 930 -285 940 -265
rect 960 -285 970 -265
rect 630 -1495 640 -325
rect 660 -1495 670 -325
rect 630 -1505 670 -1495
rect 780 -325 820 -315
rect 780 -1495 790 -325
rect 810 -1495 820 -325
rect 780 -1525 820 -1495
rect 930 -325 970 -285
rect 1230 -265 1270 -255
rect 1230 -285 1240 -265
rect 1260 -285 1270 -265
rect 930 -1495 940 -325
rect 960 -1495 970 -325
rect 930 -1505 970 -1495
rect 1080 -325 1120 -315
rect 1080 -1495 1090 -325
rect 1110 -1495 1120 -325
rect 1080 -1525 1120 -1495
rect 1230 -325 1270 -285
rect 1530 -265 1570 -255
rect 1530 -285 1540 -265
rect 1560 -285 1570 -265
rect 1230 -1495 1240 -325
rect 1260 -1495 1270 -325
rect 1230 -1505 1270 -1495
rect 1380 -325 1420 -315
rect 1380 -1495 1390 -325
rect 1410 -1495 1420 -325
rect 1380 -1525 1420 -1495
rect 1530 -325 1570 -285
rect 1830 -265 1870 -255
rect 1830 -285 1840 -265
rect 1860 -285 1870 -265
rect 1530 -1495 1540 -325
rect 1560 -1495 1570 -325
rect 1530 -1505 1570 -1495
rect 1680 -325 1720 -315
rect 1680 -1495 1690 -325
rect 1710 -1495 1720 -325
rect 1680 -1525 1720 -1495
rect 1830 -325 1870 -285
rect 2130 -265 2170 -255
rect 2130 -285 2140 -265
rect 2160 -285 2170 -265
rect 1830 -1495 1840 -325
rect 1860 -1495 1870 -325
rect 1830 -1505 1870 -1495
rect 1980 -325 2020 -315
rect 1980 -1495 1990 -325
rect 2010 -1495 2020 -325
rect 1980 -1525 2020 -1495
rect 2130 -325 2170 -285
rect 2430 -265 2470 -255
rect 2430 -285 2440 -265
rect 2460 -285 2470 -265
rect 2130 -1495 2140 -325
rect 2160 -1495 2170 -325
rect 2130 -1505 2170 -1495
rect 2280 -325 2320 -315
rect 2280 -1495 2290 -325
rect 2310 -1495 2320 -325
rect 2280 -1525 2320 -1495
rect 2430 -325 2470 -285
rect 2430 -1495 2440 -325
rect 2460 -1495 2470 -325
rect 2430 -1505 2470 -1495
rect 2580 -325 2620 -315
rect 2580 -1495 2590 -325
rect 2610 -1495 2620 -325
rect 2580 -1525 2620 -1495
rect 2660 -325 2750 -315
rect 2660 -1495 2670 -325
rect 2690 -1495 2720 -325
rect 2740 -1495 2750 -325
rect 2660 -1505 2750 -1495
rect 2860 -325 2900 -235
rect 2860 -1495 2870 -325
rect 2890 -1495 2900 -325
rect 2860 -1505 2900 -1495
rect 2940 -235 3580 -215
rect 2940 -325 2980 -235
rect 3240 -265 3280 -255
rect 3240 -285 3250 -265
rect 3270 -285 3280 -265
rect 2940 -1495 2950 -325
rect 2970 -1495 2980 -325
rect 2940 -1505 2980 -1495
rect 3090 -325 3130 -315
rect 3090 -1495 3100 -325
rect 3120 -1495 3130 -325
rect 3090 -1505 3130 -1495
rect 3240 -325 3280 -285
rect 3240 -1495 3250 -325
rect 3270 -1495 3280 -325
rect 3240 -1505 3280 -1495
rect 3390 -325 3430 -315
rect 3390 -1495 3400 -325
rect 3420 -1495 3430 -325
rect 3390 -1505 3430 -1495
rect 3540 -325 3580 -235
rect 3540 -1495 3550 -325
rect 3570 -1495 3580 -325
rect 3540 -1505 3580 -1495
rect 3620 -325 3660 -205
rect 3680 -265 3720 -255
rect 4510 -260 4550 15
rect 4660 1185 4700 1195
rect 4660 15 4670 1185
rect 4690 15 4700 1185
rect 4570 -50 4610 -40
rect 4570 -70 4580 -50
rect 4600 -55 4610 -50
rect 4660 -55 4700 15
rect 4810 1185 4850 1215
rect 4810 15 4820 1185
rect 4840 15 4850 1185
rect 4810 5 4850 15
rect 4960 1185 5000 1195
rect 4960 15 4970 1185
rect 4990 15 5000 1185
rect 4960 -55 5000 15
rect 5110 1185 5150 1195
rect 5110 15 5120 1185
rect 5140 15 5150 1185
rect 5110 -15 5150 15
rect 5260 1185 5350 1195
rect 5260 15 5270 1185
rect 5290 15 5320 1185
rect 5340 15 5350 1185
rect 5260 5 5350 15
rect 5260 -15 5300 5
rect 4600 -70 5000 -55
rect 4570 -75 5000 -70
rect 5065 -25 5150 -15
rect 5065 -45 5075 -25
rect 5095 -45 5150 -25
rect 5065 -55 5150 -45
rect 5215 -25 5300 -15
rect 5215 -45 5225 -25
rect 5245 -45 5300 -25
rect 5215 -55 5300 -45
rect 4570 -80 4610 -75
rect 5065 -105 5085 -55
rect 4570 -115 5375 -105
rect 4570 -135 4580 -115
rect 4600 -125 5375 -115
rect 4600 -135 4610 -125
rect 4570 -145 4610 -135
rect 3680 -285 3690 -265
rect 3710 -285 3720 -265
rect 3680 -295 3720 -285
rect 4220 -280 4550 -260
rect 4925 -265 5010 -255
rect 3620 -1495 3630 -325
rect 3650 -1495 3660 -325
rect 180 -1545 2620 -1525
rect 3620 -1525 3660 -1495
rect 3770 -325 3810 -315
rect 3770 -1495 3780 -325
rect 3800 -1495 3810 -325
rect 3770 -1505 3810 -1495
rect 3920 -325 3960 -315
rect 3920 -1495 3930 -325
rect 3950 -1495 3960 -325
rect 3920 -1505 3960 -1495
rect 4070 -325 4110 -315
rect 4070 -1495 4080 -325
rect 4100 -1495 4110 -325
rect 4070 -1505 4110 -1495
rect 4220 -325 4260 -280
rect 4925 -285 4935 -265
rect 4955 -285 5010 -265
rect 4925 -295 5010 -285
rect 4970 -315 5010 -295
rect 4220 -1495 4230 -325
rect 4250 -1495 4260 -325
rect 4220 -1505 4260 -1495
rect 4370 -325 4410 -315
rect 4370 -1495 4380 -325
rect 4400 -1495 4410 -325
rect 4370 -1505 4410 -1495
rect 4520 -325 4560 -315
rect 4520 -1495 4530 -325
rect 4550 -1495 4560 -325
rect 4520 -1505 4560 -1495
rect 4670 -325 4710 -315
rect 4670 -1495 4680 -325
rect 4700 -1495 4710 -325
rect 4670 -1505 4710 -1495
rect 4820 -325 4860 -315
rect 4820 -1495 4830 -325
rect 4850 -1495 4860 -325
rect 4820 -1525 4860 -1495
rect 4970 -325 5060 -315
rect 4970 -1495 4980 -325
rect 5000 -1495 5030 -325
rect 5050 -1495 5060 -325
rect 4970 -1505 5060 -1495
rect 3620 -1545 4860 -1525
<< viali >>
rect -190 15 -170 1185
rect 110 15 130 1185
rect 410 15 430 1185
rect 790 15 810 1185
rect 940 15 960 1185
rect 1090 15 1110 1185
rect -190 -1495 -170 -325
rect 110 -1495 130 -325
rect 2220 15 2240 1185
rect 2320 15 2340 1185
rect 4120 15 4140 1185
rect 4220 15 4240 1185
rect 2720 -1495 2740 -325
rect 3250 -285 3270 -265
rect 3100 -1495 3120 -325
rect 3400 -1495 3420 -325
rect 5270 15 5290 1185
rect 3690 -285 3710 -265
rect 3930 -1495 3950 -325
rect 4530 -1495 4550 -325
rect 4980 -1495 5000 -325
<< metal1 >>
rect -200 1190 -160 1195
rect -200 10 -195 1190
rect -165 10 -160 1190
rect -200 5 -160 10
rect 100 1190 140 1195
rect 100 10 105 1190
rect 135 10 140 1190
rect 100 5 140 10
rect 400 1190 440 1195
rect 400 10 405 1190
rect 435 10 440 1190
rect 400 5 440 10
rect 780 1190 820 1195
rect 780 10 785 1190
rect 815 10 820 1190
rect 780 5 820 10
rect 930 1185 970 1195
rect 930 15 940 1185
rect 960 15 970 1185
rect 930 -135 970 15
rect 1080 1190 1120 1195
rect 1080 10 1085 1190
rect 1115 10 1120 1190
rect 1080 5 1120 10
rect 2210 1190 2250 1195
rect 2210 10 2215 1190
rect 2245 10 2250 1190
rect 2210 5 2250 10
rect 2310 1190 2350 1195
rect 2310 10 2315 1190
rect 2345 10 2350 1190
rect 2310 5 2350 10
rect 4110 1190 4150 1195
rect 4110 10 4115 1190
rect 4145 10 4150 1190
rect 4110 5 4150 10
rect 4210 1190 4250 1195
rect 4210 10 4215 1190
rect 4245 10 4250 1190
rect 4210 5 4250 10
rect 5260 1190 5300 1195
rect 5260 10 5265 1190
rect 5295 10 5300 1190
rect 5260 5 5300 10
rect 930 -175 5375 -135
rect 3240 -265 3280 -175
rect 3240 -285 3250 -265
rect 3270 -285 3280 -265
rect 3240 -295 3280 -285
rect 3680 -265 3720 -175
rect 3680 -285 3690 -265
rect 3710 -285 3720 -265
rect 3680 -295 3720 -285
rect -200 -320 -160 -315
rect -200 -1500 -195 -320
rect -165 -1500 -160 -320
rect -200 -1505 -160 -1500
rect 100 -320 140 -315
rect 100 -1500 105 -320
rect 135 -1500 140 -320
rect 100 -1505 140 -1500
rect 2710 -320 2750 -315
rect 2710 -1500 2715 -320
rect 2745 -1500 2750 -320
rect 2710 -1505 2750 -1500
rect 3090 -320 3130 -315
rect 3090 -1500 3095 -320
rect 3125 -1500 3130 -320
rect 3090 -1505 3130 -1500
rect 3390 -320 3430 -315
rect 3390 -1500 3395 -320
rect 3425 -1500 3430 -320
rect 3390 -1505 3430 -1500
rect 3920 -320 3960 -315
rect 3920 -1500 3925 -320
rect 3955 -1500 3960 -320
rect 3920 -1505 3960 -1500
rect 4520 -320 4560 -315
rect 4520 -1500 4525 -320
rect 4555 -1500 4560 -320
rect 4520 -1505 4560 -1500
rect 4970 -320 5010 -315
rect 4970 -1500 4975 -320
rect 5005 -1500 5010 -320
rect 4970 -1505 5010 -1500
<< via1 >>
rect -195 1185 -165 1190
rect -195 15 -190 1185
rect -190 15 -170 1185
rect -170 15 -165 1185
rect -195 10 -165 15
rect 105 1185 135 1190
rect 105 15 110 1185
rect 110 15 130 1185
rect 130 15 135 1185
rect 105 10 135 15
rect 405 1185 435 1190
rect 405 15 410 1185
rect 410 15 430 1185
rect 430 15 435 1185
rect 405 10 435 15
rect 785 1185 815 1190
rect 785 15 790 1185
rect 790 15 810 1185
rect 810 15 815 1185
rect 785 10 815 15
rect 1085 1185 1115 1190
rect 1085 15 1090 1185
rect 1090 15 1110 1185
rect 1110 15 1115 1185
rect 1085 10 1115 15
rect 2215 1185 2245 1190
rect 2215 15 2220 1185
rect 2220 15 2240 1185
rect 2240 15 2245 1185
rect 2215 10 2245 15
rect 2315 1185 2345 1190
rect 2315 15 2320 1185
rect 2320 15 2340 1185
rect 2340 15 2345 1185
rect 2315 10 2345 15
rect 4115 1185 4145 1190
rect 4115 15 4120 1185
rect 4120 15 4140 1185
rect 4140 15 4145 1185
rect 4115 10 4145 15
rect 4215 1185 4245 1190
rect 4215 15 4220 1185
rect 4220 15 4240 1185
rect 4240 15 4245 1185
rect 4215 10 4245 15
rect 5265 1185 5295 1190
rect 5265 15 5270 1185
rect 5270 15 5290 1185
rect 5290 15 5295 1185
rect 5265 10 5295 15
rect -195 -325 -165 -320
rect -195 -1495 -190 -325
rect -190 -1495 -170 -325
rect -170 -1495 -165 -325
rect -195 -1500 -165 -1495
rect 105 -325 135 -320
rect 105 -1495 110 -325
rect 110 -1495 130 -325
rect 130 -1495 135 -325
rect 105 -1500 135 -1495
rect 2715 -325 2745 -320
rect 2715 -1495 2720 -325
rect 2720 -1495 2740 -325
rect 2740 -1495 2745 -325
rect 2715 -1500 2745 -1495
rect 3095 -325 3125 -320
rect 3095 -1495 3100 -325
rect 3100 -1495 3120 -325
rect 3120 -1495 3125 -325
rect 3095 -1500 3125 -1495
rect 3395 -325 3425 -320
rect 3395 -1495 3400 -325
rect 3400 -1495 3420 -325
rect 3420 -1495 3425 -325
rect 3395 -1500 3425 -1495
rect 3925 -325 3955 -320
rect 3925 -1495 3930 -325
rect 3930 -1495 3950 -325
rect 3950 -1495 3955 -325
rect 3925 -1500 3955 -1495
rect 4525 -325 4555 -320
rect 4525 -1495 4530 -325
rect 4530 -1495 4550 -325
rect 4550 -1495 4555 -325
rect 4525 -1500 4555 -1495
rect 4975 -325 5005 -320
rect 4975 -1495 4980 -325
rect 4980 -1495 5000 -325
rect 5000 -1495 5005 -325
rect 4975 -1500 5005 -1495
<< metal2 >>
rect -255 1190 5355 1195
rect -255 10 -195 1190
rect -165 10 105 1190
rect 135 10 405 1190
rect 435 10 785 1190
rect 815 10 1085 1190
rect 1115 10 2215 1190
rect 2245 10 2315 1190
rect 2345 10 4115 1190
rect 4145 10 4215 1190
rect 4245 10 5265 1190
rect 5295 10 5355 1190
rect -255 5 5355 10
rect -255 -320 5065 -315
rect -255 -1500 -195 -320
rect -165 -1500 105 -320
rect 135 -1500 2715 -320
rect 2745 -1500 3095 -320
rect 3125 -1500 3395 -320
rect 3425 -1500 3925 -320
rect 3955 -1500 4525 -320
rect 4555 -1500 4975 -320
rect 5005 -1500 5065 -320
rect -255 -1505 5065 -1500
<< labels >>
rlabel metal2 -255 605 -255 605 7 VP
rlabel metal2 -255 -915 -255 -915 7 VN
rlabel metal1 5375 -155 5375 -155 3 VBN
rlabel locali 5375 -115 5375 -115 3 VIN
rlabel locali 3230 1255 3230 1255 1 VOUT
rlabel locali 1400 -1545 1400 -1545 5 ROUT
<< end >>
